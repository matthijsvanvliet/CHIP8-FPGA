library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package coraxplus is

    type t_ROM is array (0 to 697 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"12", x"08", x"A4", x"65", x"DA", x"B4", x"00", x"EE", x"00", x"E0", x"68", x"32", x"6B", x"1A", x"A4", x"B1", 
        x"D8", x"B4", x"68", x"3A", x"A4", x"B5", x"D8", x"B4", x"68", x"02", x"69", x"06", x"6A", x"0B", x"6B", x"01", 
        x"65", x"2A", x"66", x"2B", x"A4", x"75", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", x"A4", x"65", x"36", x"2B", 
        x"A4", x"61", x"DA", x"B4", x"6B", x"06", x"A4", x"79", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", x"A4", x"61", 
        x"45", x"2A", x"A4", x"65", x"DA", x"B4", x"6B", x"0B", x"A4", x"7D", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", 
        x"A4", x"61", x"55", x"60", x"A4", x"65", x"DA", x"B4", x"6B", x"10", x"A4", x"85", x"D8", x"B4", x"A4", x"AD", 
        x"D9", x"B4", x"A4", x"61", x"76", x"FF", x"46", x"2A", x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"8D", 
        x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", x"A4", x"61", x"95", x"60", x"A4", x"65", x"DA", x"B4", x"7B", x"05", 
        x"A4", x"6D", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", x"A4", x"65", x"12", x"8E", x"A4", x"61", x"DA", x"B4", 
        x"68", x"12", x"69", x"16", x"6A", x"1B", x"6B", x"01", x"A4", x"71", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", 
        x"22", x"02", x"7B", x"05", x"A4", x"69", x"D8", x"B4", x"A4", x"A1", x"D9", x"B4", x"A4", x"65", x"DA", x"B4", 
        x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"69", x"D9", x"B4", x"A4", x"61", x"65", x"2A", x"67", x"00", 
        x"87", x"50", x"47", x"2A", x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"6D", 
        x"D9", x"B4", x"A4", x"61", x"66", x"0B", x"67", x"2A", x"87", x"61", x"47", x"2B", x"A4", x"65", x"DA", x"B4", 
        x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"71", x"D9", x"B4", x"A4", x"61", x"66", x"78", x"67", x"1F", 
        x"87", x"62", x"47", x"18", x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"75", 
        x"D9", x"B4", x"A4", x"61", x"66", x"78", x"67", x"1F", x"87", x"63", x"47", x"67", x"A4", x"65", x"DA", x"B4", 
        x"68", x"22", x"69", x"26", x"6A", x"2B", x"6B", x"01", x"A4", x"89", x"D8", x"B4", x"A4", x"79", x"D9", x"B4", 
        x"A4", x"61", x"66", x"8C", x"67", x"8C", x"87", x"64", x"47", x"18", x"A4", x"65", x"DA", x"B4", x"7B", x"05", 
        x"A4", x"89", x"D8", x"B4", x"A4", x"7D", x"D9", x"B4", x"A4", x"61", x"66", x"8C", x"67", x"78", x"87", x"65", 
        x"47", x"EC", x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"85", x"D9", x"B4", 
        x"A4", x"61", x"66", x"78", x"67", x"8C", x"87", x"67", x"47", x"EC", x"A4", x"65", x"DA", x"B4", x"7B", x"05", 
        x"A4", x"89", x"D8", x"B4", x"A4", x"81", x"D9", x"B4", x"A4", x"61", x"66", x"0F", x"86", x"66", x"46", x"07", 
        x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"89", x"D8", x"B4", x"A4", x"A1", x"D9", x"B4", x"A4", x"61", 
        x"66", x"E0", x"86", x"6E", x"46", x"C0", x"A4", x"65", x"DA", x"B4", x"7B", x"05", x"A4", x"A5", x"D8", x"B4", 
        x"A4", x"81", x"D9", x"B4", x"A4", x"5E", x"F1", x"65", x"A4", x"65", x"30", x"AA", x"A4", x"61", x"31", x"55", 
        x"A4", x"61", x"DA", x"B4", x"68", x"32", x"69", x"36", x"6A", x"3B", x"6B", x"01", x"A4", x"A5", x"D8", x"B4", 
        x"A4", x"7D", x"D9", x"B4", x"A4", x"5E", x"60", x"00", x"61", x"30", x"F1", x"55", x"A4", x"5E", x"F0", x"65", 
        x"81", x"00", x"A4", x"5F", x"F0", x"65", x"A4", x"65", x"30", x"30", x"A4", x"61", x"31", x"00", x"A4", x"61", 
        x"DA", x"B4", x"7B", x"05", x"A4", x"A5", x"D8", x"B4", x"A4", x"75", x"D9", x"B4", x"A4", x"5E", x"66", x"89", 
        x"F6", x"33", x"F2", x"65", x"A4", x"65", x"30", x"01", x"A4", x"61", x"31", x"03", x"A4", x"61", x"32", x"07", 
        x"A4", x"61", x"DA", x"B4", x"7B", x"05", x"A4", x"A5", x"D8", x"B4", x"A4", x"A1", x"D9", x"B4", x"A4", x"61", 
        x"66", x"04", x"F6", x"1E", x"DA", x"B4", x"7B", x"05", x"A4", x"A9", x"D8", x"B4", x"A4", x"AD", x"D9", x"B4", 
        x"A4", x"65", x"66", x"FF", x"76", x"0A", x"36", x"09", x"A4", x"61", x"86", x"66", x"36", x"04", x"A4", x"61", 
        x"66", x"FF", x"60", x"0A", x"86", x"04", x"36", x"09", x"A4", x"61", x"86", x"66", x"36", x"04", x"A4", x"61", 
        x"66", x"FF", x"86", x"6E", x"86", x"66", x"36", x"7F", x"A4", x"61", x"86", x"66", x"86", x"6E", x"36", x"7E", 
        x"A4", x"61", x"66", x"05", x"76", x"F6", x"36", x"FB", x"A4", x"61", x"66", x"05", x"86", x"05", x"36", x"FB", 
        x"A4", x"61", x"66", x"05", x"80", x"67", x"30", x"FB", x"A4", x"61", x"DA", x"B4", x"14", x"5C", x"AA", x"55", 
        x"00", x"00", x"A0", x"40", x"A0", x"00", x"A0", x"C0", x"80", x"E0", x"A0", x"A0", x"E0", x"C0", x"40", x"40", 
        x"E0", x"E0", x"20", x"C0", x"E0", x"E0", x"60", x"20", x"E0", x"A0", x"E0", x"20", x"20", x"E0", x"C0", x"20", 
        x"C0", x"60", x"80", x"E0", x"E0", x"E0", x"20", x"40", x"40", x"E0", x"E0", x"A0", x"E0", x"E0", x"E0", x"20", 
        x"C0", x"40", x"A0", x"E0", x"A0", x"C0", x"E0", x"A0", x"E0", x"E0", x"80", x"80", x"E0", x"C0", x"A0", x"A0", 
        x"C0", x"E0", x"C0", x"80", x"E0", x"E0", x"80", x"C0", x"80", x"00", x"A0", x"A0", x"40", x"A0", x"40", x"A0", 
        x"A0", x"0A", x"AE", x"A2", x"42", x"38", x"28", x"28", x"B8"
    );

end package;

package body coraxplus is
end coraxplus;