library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package down8 is

    type t_ROM is array (0 to 2017 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"14", x"36", x"47", x"01", x"00", x"EE", x"67", x"01", x"65", x"FE", x"22", x"54", x"76", x"01", x"A4", x"EA", 
        x"F6", x"33", x"22", x"54", x"A4", x"EE", x"F2", x"65", x"6F", x"09", x"8F", x"45", x"4F", x"00", x"12", x"26", 
        x"69", x"08", x"88", x"00", x"12", x"38", x"6F", x"11", x"8F", x"45", x"4F", x"00", x"12", x"34", x"69", x"10", 
        x"88", x"10", x"12", x"38", x"69", x"18", x"88", x"20", x"A4", x"F1", x"F0", x"65", x"A4", x"E2", x"6F", x"0A", 
        x"8F", x"07", x"3F", x"00", x"A4", x"E4", x"6F", x"14", x"8F", x"07", x"3F", x"00", x"A4", x"E6", x"D8", x"92", 
        x"6C", x"01", x"00", x"EE", x"A4", x"EA", x"F2", x"65", x"68", x"31", x"69", x"1A", x"F0", x"29", x"D8", x"95", 
        x"78", x"05", x"F1", x"29", x"D8", x"95", x"78", x"05", x"F2", x"29", x"D8", x"95", x"78", x"F6", x"00", x"EE", 
        x"A4", x"F1", x"F0", x"65", x"70", x"01", x"A4", x"F1", x"F0", x"55", x"00", x"E0", x"23", x"0E", x"22", x"54", 
        x"23", x"5C", x"A4", x"F1", x"F0", x"65", x"A4", x"E2", x"6F", x"0A", x"8F", x"07", x"3F", x"00", x"A4", x"E4", 
        x"6F", x"14", x"8F", x"07", x"3F", x"00", x"A4", x"E6", x"69", x"08", x"C8", x"0F", x"78", x"0C", x"80", x"80", 
        x"D8", x"92", x"69", x"10", x"C8", x"0F", x"78", x"0C", x"81", x"80", x"D8", x"92", x"69", x"18", x"C8", x"0F", 
        x"78", x"0C", x"82", x"80", x"D8", x"92", x"64", x"00", x"A4", x"EE", x"F2", x"55", x"A4", x"E0", x"D3", x"42", 
        x"6F", x"14", x"22", x"C6", x"00", x"EE", x"FF", x"15", x"FF", x"07", x"3F", x"00", x"12", x"C8", x"00", x"EE", 
        x"75", x"01", x"45", x"01", x"67", x"00", x"00", x"EE", x"A4", x"EE", x"F2", x"65", x"40", x"00", x"00", x"EE", 
        x"3C", x"00", x"13", x"0A", x"6F", x"0A", x"FF", x"18", x"A4", x"ED", x"F0", x"65", x"8F", x"60", x"8F", x"07", 
        x"4F", x"00", x"80", x"60", x"A4", x"ED", x"F0", x"55", x"66", x"00", x"22", x"54", x"A4", x"EA", x"F6", x"33", 
        x"22", x"54", x"23", x"5C", x"7D", x"FF", x"3D", x"FF", x"23", x"5C", x"6C", x"00", x"00", x"EE", x"A4", x"F1", 
        x"F0", x"65", x"68", x"00", x"69", x"00", x"A4", x"F5", x"6F", x"0A", x"8F", x"07", x"3F", x"00", x"A5", x"05", 
        x"6F", x"14", x"8F", x"07", x"3F", x"00", x"A5", x"0D", x"D8", x"98", x"79", x"08", x"D8", x"98", x"79", x"08", 
        x"D8", x"98", x"79", x"08", x"D8", x"98", x"68", x"21", x"69", x"00", x"A4", x"FD", x"6F", x"0A", x"8F", x"07", 
        x"3F", x"00", x"A5", x"05", x"6F", x"14", x"8F", x"07", x"3F", x"00", x"A5", x"15", x"D8", x"98", x"79", x"08", 
        x"D8", x"98", x"79", x"08", x"D8", x"98", x"79", x"08", x"D8", x"98", x"00", x"EE", x"68", x"39", x"69", x"01", 
        x"FD", x"29", x"D8", x"95", x"79", x"05", x"A5", x"1D", x"D8", x"93", x"79", x"04", x"68", x"04", x"F8", x"29", 
        x"68", x"3B", x"D8", x"95", x"A4", x"E0", x"00", x"EE", x"6A", x"00", x"6B", x"00", x"6C", x"08", x"DA", x"B8", 
        x"FC", x"1E", x"8A", x"C4", x"4A", x"40", x"7B", x"08", x"4A", x"40", x"6A", x"00", x"3B", x"20", x"13", x"7E", 
        x"00", x"EE", x"6F", x"1E", x"22", x"C6", x"00", x"E0", x"A5", x"4A", x"23", x"78", x"A4", x"ED", x"F0", x"65", 
        x"A4", x"EA", x"F0", x"33", x"22", x"54", x"A4", x"F1", x"F0", x"65", x"F0", x"33", x"F2", x"65", x"68", x"01", 
        x"69", x"01", x"A5", x"2F", x"D8", x"95", x"78", x"05", x"A5", x"33", x"D8", x"95", x"78", x"05", x"A5", x"38", 
        x"D8", x"95", x"78", x"0A", x"F1", x"29", x"D8", x"95", x"78", x"05", x"69", x"03", x"A5", x"33", x"D8", x"91", 
        x"F2", x"29", x"78", x"05", x"69", x"01", x"D8", x"95", x"68", x"1A", x"69", x"1A", x"A5", x"20", x"D8", x"95", 
        x"78", x"06", x"A5", x"25", x"D8", x"95", x"78", x"06", x"A5", x"2A", x"D8", x"95", x"66", x"00", x"A4", x"EA", 
        x"F6", x"33", x"A4", x"EE", x"60", x"00", x"61", x"00", x"62", x"00", x"F2", x"55", x"A4", x"F1", x"F0", x"55", 
        x"6A", x"05", x"EA", x"A1", x"14", x"74", x"14", x"00", x"A4", x"F1", x"F0", x"65", x"30", x"00", x"14", x"14", 
        x"60", x"28", x"14", x"16", x"60", x"00", x"A4", x"F1", x"F0", x"55", x"68", x"14", x"69", x"14", x"A5", x"3D", 
        x"D8", x"95", x"A5", x"42", x"78", x"04", x"D8", x"94", x"A5", x"46", x"78", x"04", x"D8", x"94", x"78", x"03", 
        x"D8", x"94", x"A4", x"DE", x"00", x"EE", x"A6", x"4A", x"23", x"78", x"63", x"04", x"64", x"00", x"A4", x"E0", 
        x"D3", x"42", x"A4", x"DE", x"D3", x"43", x"74", x"01", x"6A", x"0F", x"EA", x"A1", x"24", x"08", x"6A", x"05", 
        x"EA", x"A1", x"14", x"5A", x"6F", x"03", x"22", x"C6", x"14", x"44", x"00", x"E0", x"A7", x"4A", x"23", x"78", 
        x"A4", x"E8", x"63", x"2D", x"64", x"17", x"D3", x"42", x"6A", x"05", x"EA", x"A1", x"14", x"74", x"6F", x"14", 
        x"22", x"C6", x"14", x"66", x"00", x"E0", x"23", x"0E", x"63", x"13", x"64", x"00", x"6C", x"00", x"65", x"01", 
        x"6D", x"04", x"22", x"54", x"23", x"5C", x"A4", x"E0", x"D3", x"42", x"D3", x"42", x"6A", x"09", x"EA", x"A1", 
        x"73", x"01", x"6A", x"07", x"EA", x"A1", x"73", x"FF", x"43", x"07", x"73", x"01", x"43", x"20", x"73", x"FF", 
        x"84", x"54", x"35", x"02", x"75", x"01", x"6A", x"05", x"EA", x"9E", x"14", x"B0", x"67", x"01", x"14", x"B2", 
        x"67", x"00", x"D3", x"42", x"4F", x"01", x"22", x"02", x"44", x"0A", x"22", x"D8", x"44", x"12", x"22", x"D8", 
        x"44", x"1A", x"22", x"D8", x"A4", x"E0", x"6F", x"1F", x"8F", x"47", x"3F", x"00", x"22", x"70", x"4D", x"FF", 
        x"13", x"92", x"FF", x"07", x"3F", x"00", x"14", x"D2", x"6F", x"03", x"FF", x"15", x"14", x"8A", x"C0", x"00", 
        x"C0", x"C0", x"F0", x"60", x"E0", x"40", x"40", x"40", x"41", x"22", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"1E", x"AB", x"55", x"01", x"2B", x"01", x"55", x"01", x"70", x"AA", x"D4", 
        x"80", x"AA", x"80", x"D4", x"80", x"FE", x"01", x"7F", x"80", x"FE", x"01", x"7F", x"80", x"15", x"09", x"01", 
        x"85", x"41", x"81", x"01", x"09", x"82", x"85", x"82", x"80", x"90", x"A8", x"91", x"80", x"04", x"38", x"40", 
        x"50", x"A8", x"A8", x"A8", x"88", x"70", x"48", x"88", x"F8", x"88", x"80", x"58", x"20", x"50", x"C8", x"80", 
        x"80", x"80", x"80", x"F0", x"80", x"E0", x"80", x"F0", x"90", x"90", x"A0", x"60", x"40", x"C0", x"A0", x"C0", 
        x"A0", x"C0", x"E0", x"A0", x"A0", x"E0", x"40", x"80", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"0A", x"0A", x"0A", x"0A", x"0A", x"0A", 
        x"0A", x"F2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"51", x"00", x"04", 
        x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"FF", x"00", x"00", x"00", x"00", 
        x"00", x"08", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"8F", x"00", x"FF", x"00", x"00", x"00", x"00", 
        x"00", x"22", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"F8", x"00", x"00", x"08", x"08", 
        x"08", x"79", x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"C1", x"01", x"02", x"00", x"00", x"00", x"00", 
        x"00", x"E3", x"40", x"80", x"00", x"00", x"40", x"40", x"40", x"C0", x"08", x"0D", x"05", x"05", x"02", x"02", 
        x"04", x"1C", x"99", x"10", x"10", x"19", x"0F", x"00", x"00", x"00", x"A2", x"A2", x"A2", x"A6", x"1E", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"88", x"88", x"88", x"98", x"69", x"00", 
        x"00", x"00", x"42", x"43", x"42", x"43", x"F1", x"00", x"00", x"00", x"14", x"F4", x"04", x"04", x"F3", x"00", 
        x"00", x"00", x"40", x"40", x"40", x"C6", x"46", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"20", x"02", x"00", x"1C", x"22", x"41", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"7F", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"61", x"81", x"A0", x"81", x"A0", x"81", 
        x"A0", x"81", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"30", x"30", x"30", 
        x"30", x"30", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"1E", x"7F", 
        x"61", x"61", x"FE", x"01", x"01", x"01", x"01", x"01", x"81", x"81", x"A0", x"81", x"A0", x"81", x"A0", x"81", 
        x"A0", x"81", x"03", x"07", x"0E", x"0C", x"0C", x"0E", x"07", x"03", x"F1", x"F3", x"36", x"36", x"36", x"36", 
        x"F3", x"F1", x"C6", x"E6", x"36", x"36", x"36", x"36", x"E3", x"C3", x"66", x"66", x"66", x"F6", x"D6", x"D6", 
        x"9C", x"9C", x"DC", x"FE", x"E6", x"C6", x"C6", x"C6", x"C6", x"C6", x"7F", x"3F", x"73", x"61", x"61", x"61", 
        x"7F", x"1E", x"01", x"01", x"81", x"81", x"81", x"81", x"01", x"01", x"A0", x"81", x"A0", x"81", x"A0", x"81", 
        x"A0", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"03", x"02", x"02", x"00", x"00", x"00", x"00", x"00", x"01", 
        x"44", x"54", x"01", x"01", x"01", x"01", x"01", x"81", x"81", x"81", x"A0", x"81", x"A0", x"81", x"A0", x"81", 
        x"A0", x"61", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"FF", x"02", x"02", x"03", x"00", x"00", x"00", x"00", x"FF", x"54", x"28", x"01", x"00", x"00", x"00", 
        x"00", x"FF", x"81", x"81", x"81", x"01", x"01", x"01", x"01", x"FE", x"7F", x"80", x"80", x"80", x"80", x"8F", 
        x"90", x"93", x"FF", x"00", x"00", x"00", x"00", x"00", x"F0", x"8F", x"FF", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"87", x"FF", x"00", x"00", x"00", x"00", x"03", x"3C", x"C7", x"FF", x"00", x"00", x"00", x"01", x"C1", 
        x"21", x"21", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"24", x"FF", x"00", x"0F", x"F8", x"00", x"00", 
        x"00", x"E7", x"FE", x"01", x"E1", x"11", x"11", x"11", x"11", x"11", x"94", x"94", x"94", x"94", x"94", x"94", 
        x"94", x"94", x"00", x"00", x"06", x"09", x"09", x"0F", x"09", x"00", x"48", x"30", x"03", x"02", x"32", x"02", 
        x"03", x"30", x"00", x"00", x"80", x"40", x"40", x"40", x"80", x"00", x"A1", x"A1", x"A1", x"A1", x"A1", x"A1", 
        x"A1", x"A1", x"24", x"3C", x"24", x"24", x"00", x"00", x"00", x"00", x"42", x"42", x"42", x"E2", x"00", x"00", 
        x"00", x"40", x"11", x"11", x"11", x"11", x"11", x"11", x"11", x"11", x"94", x"94", x"94", x"94", x"94", x"94", 
        x"94", x"94", x"00", x"10", x"20", x"7F", x"20", x"10", x"00", x"00", x"00", x"00", x"30", x"03", x"00", x"30", 
        x"00", x"00", x"00", x"20", x"10", x"F8", x"10", x"20", x"00", x"00", x"A1", x"A1", x"A1", x"A1", x"A1", x"A1", 
        x"A1", x"A1", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"03", x"40", x"50", x"E0", x"40", x"00", x"00", 
        x"00", x"F0", x"11", x"11", x"11", x"11", x"11", x"11", x"31", x"11", x"94", x"94", x"8B", x"87", x"80", x"80", 
        x"80", x"7F", x"00", x"78", x"C7", x"F0", x"0F", x"00", x"00", x"FF", x"30", x"00", x"87", x"FC", x"FF", x"00", 
        x"00", x"FF", x"00", x"78", x"8F", x"7F", x"80", x"00", x"00", x"FF", x"A1", x"A1", x"C1", x"00", x"00", x"00", 
        x"00", x"FF", x"01", x"00", x"80", x"83", x"BC", x"60", x"00", x"FF", x"E0", x"00", x"00", x"FF", x"00", x"00", 
        x"00", x"FF", x"11", x"11", x"51", x"11", x"F1", x"01", x"01", x"FE"
    );

end package;

package body down8 is
end down8;