library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package danm8ku is

    type t_ROM is array (0 to 2017 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"14", x"E2", x"E0", x"00", x"80", x"79", x"00", x"60", x"0C", x"0C", x"3E", x"0C", x"9B", x"FD", x"20", x"63", 
        x"1C", x"0C", x"3E", x"0C", x"FB", x"CD", x"70", x"E7", x"1C", x"1E", x"23", x"0C", x"F3", x"FD", x"F8", x"CF", 
        x"1E", x"1F", x"21", x"0C", x"C3", x"FD", x"D8", x"CD", x"1E", x"9B", x"21", x"1C", x"E3", x"CD", x"DD", x"DD", 
        x"9E", x"BF", x"21", x"98", x"F3", x"8D", x"CD", x"D9", x"9F", x"3F", x"23", x"F8", x"F9", x"9D", x"CD", x"D9", 
        x"DB", x"71", x"3F", x"F0", x"98", x"F9", x"CD", x"D9", x"D9", x"60", x"3C", x"00", x"00", x"F8", x"00", x"00", 
        x"00", x"00", x"00", x"1E", x"10", x"10", x"10", x"1E", x"10", x"10", x"10", x"EA", x"AA", x"AA", x"AA", x"EE", 
        x"EA", x"8A", x"8E", x"8A", x"EA", x"AE", x"A8", x"4C", x"48", x"4E", x"E4", x"84", x"E4", x"20", x"E4", x"FF", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A0", x"A0", x"00", x"00", x"50", x"50", x"00", x"00", x"60", 
        x"60", x"00", x"60", x"00", x"60", x"00", x"C0", x"A0", x"60", x"00", x"30", x"50", x"60", x"00", x"00", x"05", 
        x"0F", x"00", x"00", x"60", x"00", x"60", x"00", x"60", x"A0", x"C0", x"00", x"60", x"50", x"30", x"00", x"60", 
        x"60", x"00", x"00", x"C0", x"C0", x"00", x"00", x"30", x"30", x"00", x"C0", x"60", x"C0", x"00", x"60", x"60", 
        x"00", x"00", x"C0", x"C0", x"00", x"00", x"30", x"30", x"00", x"00", x"A0", x"40", x"A0", x"00", x"00", x"00", 
        x"60", x"60", x"00", x"00", x"C0", x"C0", x"00", x"00", x"30", x"30", x"00", x"E0", x"6A", x"38", x"6B", x"0B", 
        x"A2", x"03", x"DA", x"B1", x"F0", x"65", x"7A", x"F8", x"4A", x"F8", x"7B", x"01", x"4A", x"F8", x"6A", x"38", 
        x"3B", x"15", x"12", x"D2", x"64", x"05", x"E4", x"A1", x"00", x"EE", x"64", x"07", x"E4", x"A1", x"00", x"EE", 
        x"64", x"08", x"E4", x"A1", x"00", x"EE", x"64", x"09", x"E4", x"A1", x"00", x"EE", x"A2", x"02", x"60", x"00", 
        x"C1", x"1F", x"71", x"F6", x"6F", x"0B", x"8F", x"17", x"4F", x"00", x"12", x"E4", x"71", x"0A", x"62", x"3C", 
        x"40", x"20", x"12", x"E4", x"D0", x"12", x"D2", x"12", x"3F", x"01", x"12", x"E4", x"70", x"04", x"72", x"FC", 
        x"13", x"10", x"00", x"E0", x"63", x"1F", x"65", x"3F", x"A2", x"65", x"60", x"1A", x"61", x"0E", x"D0", x"15", 
        x"70", x"08", x"A2", x"6A", x"D0", x"15", x"A0", x"00", x"60", x"03", x"61", x"01", x"62", x"20", x"66", x"20", 
        x"64", x"20", x"82", x"04", x"86", x"05", x"84", x"15", x"87", x"20", x"8B", x"10", x"23", x"66", x"87", x"60", 
        x"23", x"66", x"8B", x"40", x"23", x"66", x"87", x"20", x"23", x"66", x"70", x"01", x"71", x"01", x"40", x"20", 
        x"70", x"01", x"80", x"52", x"13", x"3C", x"8B", x"32", x"87", x"52", x"6C", x"00", x"6F", x"15", x"8F", x"77", 
        x"4F", x"00", x"7C", x"01", x"6F", x"29", x"8F", x"75", x"4F", x"00", x"7C", x"01", x"6F", x"0A", x"8F", x"B7", 
        x"4F", x"00", x"7C", x"01", x"6F", x"13", x"8F", x"B5", x"4F", x"00", x"7C", x"01", x"6F", x"00", x"8F", x"C5", 
        x"4F", x"00", x"D7", x"B4", x"00", x"EE", x"00", x"E0", x"A2", x"5B", x"60", x"19", x"61", x"0D", x"D0", x"15", 
        x"A2", x"60", x"70", x"08", x"D0", x"15", x"F0", x"0A", x"F0", x"0A", x"00", x"EE", x"60", x"FF", x"24", x"20", 
        x"A2", x"9E", x"83", x"3E", x"83", x"3E", x"F3", x"1E", x"D4", x"54", x"00", x"EE", x"8C", x"00", x"80", x"0E", 
        x"8A", x"F0", x"86", x"04", x"80", x"C0", x"8A", x"F2", x"88", x"F0", x"88", x"A5", x"88", x"A5", x"84", x"84", 
        x"8C", x"10", x"81", x"1E", x"8A", x"F0", x"87", x"14", x"81", x"C0", x"8A", x"F2", x"8D", x"F0", x"8D", x"A5", 
        x"8D", x"A5", x"85", x"D4", x"6F", x"FA", x"8F", x"07", x"3F", x"00", x"13", x"F2", x"80", x"24", x"3F", x"00", 
        x"80", x"25", x"83", x"80", x"6F", x"01", x"8F", x"85", x"4F", x"00", x"63", x"02", x"6F", x"01", x"8F", x"D5", 
        x"4F", x"00", x"6D", x"02", x"8D", x"DE", x"8D", x"DE", x"83", x"D1", x"6F", x"3E", x"8F", x"45", x"3F", x"00", 
        x"14", x"16", x"23", x"AC", x"14", x"1E", x"6F", x"1D", x"8F", x"55", x"4F", x"00", x"23", x"AC", x"00", x"EE", 
        x"AB", x"B8", x"FB", x"1E", x"F7", x"55", x"00", x"EE", x"6B", x"00", x"AB", x"B8", x"FB", x"1E", x"F7", x"65", 
        x"40", x"FF", x"14", x"3E", x"A2", x"72", x"83", x"3E", x"83", x"3E", x"F3", x"1E", x"D4", x"54", x"7B", x"08", 
        x"3B", x"00", x"14", x"2A", x"00", x"EE", x"6B", x"00", x"AB", x"B8", x"FB", x"1E", x"F7", x"65", x"30", x"FF", 
        x"23", x"BC", x"30", x"FF", x"24", x"20", x"7B", x"08", x"3B", x"00", x"14", x"48", x"00", x"EE", x"AB", x"54", 
        x"F7", x"55", x"A2", x"8E", x"F0", x"65", x"AB", x"B8", x"F0", x"1E", x"F7", x"65", x"68", x"00", x"30", x"FF", 
        x"14", x"80", x"A2", x"8E", x"F0", x"65", x"8A", x"00", x"70", x"08", x"A2", x"8E", x"F0", x"55", x"68", x"01", 
        x"AB", x"54", x"F7", x"65", x"63", x"00", x"AB", x"B8", x"FA", x"1E", x"00", x"EE", x"FF", x"07", x"3F", x"00", 
        x"14", x"8C", x"6F", x"01", x"FF", x"15", x"00", x"EE", x"A2", x"8F", x"F1", x"65", x"83", x"16", x"82", x"06", 
        x"A2", x"AA", x"D2", x"33", x"62", x"05", x"E2", x"9E", x"14", x"B0", x"71", x"FF", x"41", x"01", x"61", x"02", 
        x"62", x"07", x"E2", x"9E", x"14", x"BC", x"70", x"FF", x"40", x"01", x"60", x"02", x"62", x"09", x"E2", x"9E", 
        x"14", x"C8", x"70", x"01", x"40", x"23", x"60", x"22", x"62", x"08", x"E2", x"9E", x"14", x"D4", x"71", x"01", 
        x"41", x"3A", x"61", x"39", x"A2", x"8F", x"F1", x"55", x"83", x"16", x"82", x"06", x"A2", x"AA", x"D2", x"33", 
        x"00", x"EE", x"22", x"CA", x"69", x"00", x"60", x"00", x"A2", x"AD", x"F0", x"55", x"6B", x"00", x"A2", x"6F", 
        x"F7", x"65", x"AB", x"B8", x"F7", x"55", x"7B", x"01", x"3B", x"20", x"14", x"F4", x"00", x"E0", x"A2", x"53", 
        x"60", x"39", x"61", x"00", x"D0", x"18", x"71", x"08", x"6F", x"20", x"8F", x"17", x"4F", x"00", x"15", x"04", 
        x"A2", x"8F", x"F1", x"65", x"83", x"16", x"82", x"06", x"A2", x"AA", x"D2", x"33", x"24", x"28", x"24", x"98", 
        x"4F", x"01", x"15", x"34", x"24", x"46", x"8D", x"90", x"25", x"5C", x"4D", x"FF", x"25", x"38", x"79", x"01", 
        x"24", x"8C", x"15", x"1C", x"23", x"96", x"14", x"E2", x"A2", x"AD", x"F0", x"65", x"70", x"01", x"A2", x"AD", 
        x"F0", x"55", x"62", x"3D", x"61", x"01", x"80", x"06", x"3F", x"00", x"15", x"5A", x"40", x"01", x"15", x"56", 
        x"71", x"04", x"70", x"FF", x"15", x"4C", x"A2", x"BA", x"D2", x"13", x"00", x"EE", x"A2", x"AD", x"F0", x"65", 
        x"6F", x"01", x"80", x"F2", x"30", x"01", x"15", x"6E", x"4D", x"8C", x"69", x"FE", x"15", x"74", x"A2", x"AD", 
        x"F0", x"65", x"B7", x"15", x"00", x"EE", x"F7", x"55", x"A2", x"7E", x"D4", x"54", x"00", x"EE", x"60", x"07", 
        x"80", x"D2", x"30", x"07", x"15", x"96", x"CC", x"1F", x"24", x"5E", x"62", x"02", x"C0", x"3F", x"70", x"AA", 
        x"64", x"37", x"85", x"C0", x"25", x"76", x"15", x"74", x"60", x"03", x"80", x"D2", x"30", x"03", x"15", x"CC", 
        x"CC", x"1F", x"24", x"5E", x"38", x"01", x"15", x"B6", x"C0", x"7F", x"70", x"7F", x"64", x"39", x"85", x"C0", 
        x"61", x"23", x"62", x"00", x"25", x"76", x"CC", x"1F", x"24", x"5E", x"38", x"01", x"15", x"CC", x"C0", x"7F", 
        x"70", x"7F", x"64", x"39", x"85", x"C0", x"61", x"9B", x"62", x"00", x"25", x"76", x"15", x"74", x"00", x"00", 
        x"00", x"CE", x"32", x"D2", x"2E", x"D6", x"2A", x"DA", x"26", x"DE", x"22", x"E2", x"1E", x"E6", x"1A", x"EA", 
        x"16", x"EE", x"12", x"F2", x"0E", x"F6", x"0A", x"FA", x"06", x"FE", x"02", x"FA", x"82", x"F6", x"86", x"F2", 
        x"8A", x"EE", x"8E", x"EA", x"92", x"E6", x"96", x"E2", x"9A", x"DE", x"9E", x"DA", x"A2", x"D6", x"A6", x"D2", 
        x"AA", x"CE", x"AE", x"A5", x"CE", x"FD", x"33", x"A5", x"CE", x"F2", x"65", x"32", x"00", x"16", x"25", x"40", 
        x"01", x"71", x"0A", x"40", x"02", x"71", x"14", x"81", x"1E", x"F1", x"1E", x"F1", x"65", x"24", x"5E", x"64", 
        x"3C", x"65", x"10", x"25", x"76", x"15", x"74", x"60", x"0F", x"80", x"D2", x"30", x"0F", x"16", x"55", x"CC", 
        x"1F", x"64", x"3C", x"85", x"C0", x"60", x"96", x"61", x"00", x"24", x"5E", x"62", x"08", x"25", x"76", x"24", 
        x"5E", x"62", x"04", x"25", x"76", x"64", x"2D", x"60", x"4B", x"24", x"5E", x"61", x"87", x"25", x"76", x"24", 
        x"5E", x"61", x"0A", x"25", x"76", x"15", x"74", x"CC", x"1F", x"24", x"5E", x"64", x"32", x"85", x"C0", x"60", 
        x"E6", x"61", x"00", x"25", x"76", x"24", x"5E", x"64", x"36", x"25", x"76", x"24", x"5E", x"64", x"3A", x"25", 
        x"76", x"00", x"EE", x"60", x"1F", x"80", x"D2", x"30", x"1F", x"16", x"91", x"CC", x"1F", x"24", x"5E", x"64", 
        x"23", x"85", x"C0", x"60", x"42", x"61", x"0C", x"62", x"02", x"25", x"76", x"24", x"5E", x"61", x"82", x"25", 
        x"76", x"4D", x"40", x"26", x"57", x"4D", x"80", x"26", x"57", x"4D", x"C0", x"26", x"57", x"15", x"74", x"60", 
        x"07", x"80", x"D2", x"30", x"07", x"16", x"C3", x"60", x"20", x"80", x"D2", x"40", x"00", x"16", x"B5", x"65", 
        x"1C", x"61", x"A0", x"16", x"B9", x"65", x"00", x"61", x"1E", x"C4", x"1F", x"74", x"1F", x"60", x"BE", x"24", 
        x"5E", x"25", x"76", x"15", x"74", x"60", x"07", x"80", x"D2", x"30", x"07", x"16", x"E7", x"60", x"10", x"80", 
        x"D2", x"65", x"1C", x"61", x"A0", x"30", x"00", x"16", x"DD", x"65", x"00", x"61", x"1E", x"60", x"00", x"62", 
        x"00", x"C4", x"1F", x"24", x"5E", x"25", x"76", x"15", x"74", x"60", x"0F", x"80", x"D2", x"30", x"0F", x"17", 
        x"0F", x"85", x"D6", x"85", x"56", x"85", x"56", x"64", x"32", x"60", x"5F", x"61", x"00", x"62", x"05", x"24", 
        x"5E", x"25", x"76", x"61", x"14", x"24", x"5E", x"25", x"76", x"61", x"94", x"24", x"5E", x"25", x"76", x"15", 
        x"74", x"23", x"22", x"14", x"E2", x"15", x"7E", x"15", x"98", x"16", x"03", x"16", x"27", x"16", x"73", x"16", 
        x"9F", x"16", x"C5", x"16", x"E9", x"17", x"11"
    );

end package;

package body danm8ku is
end danm8ku;