library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package octojam9title is

    type t_ROM is array (0 to 690 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"60", x"10", x"62", x"0B", x"A3", x"F6", x"D0", x"1B", x"F2", x"1E", x"81", x"24", x"41", x"21", x"70", x"08", 
        x"41", x"21", x"61", x"00", x"30", x"30", x"12", x"06", x"23", x"E6", x"62", x"08", x"60", x"12", x"61", x"02", 
        x"D0", x"18", x"23", x"EA", x"F2", x"1E", x"60", x"1C", x"61", x"02", x"D0", x"18", x"23", x"EA", x"F2", x"1E", 
        x"60", x"26", x"61", x"02", x"D0", x"18", x"23", x"EA", x"F2", x"1E", x"60", x"26", x"61", x"0C", x"D0", x"18", 
        x"23", x"EA", x"F2", x"1E", x"60", x"26", x"61", x"16", x"D0", x"18", x"23", x"EA", x"F2", x"1E", x"60", x"1C", 
        x"61", x"16", x"D0", x"18", x"23", x"EA", x"F2", x"1E", x"60", x"12", x"61", x"16", x"D0", x"18", x"23", x"EA", 
        x"F2", x"1E", x"23", x"E6", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"12", x"61", x"02", x"D0", x"18", x"71", x"02", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"06", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"02", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"1C", x"61", x"02", x"D0", x"18", x"70", x"FE", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"FA", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"FE", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"26", x"61", x"02", x"D0", x"18", x"70", x"FE", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"FA", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"FE", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"26", x"61", x"0C", x"D0", x"18", x"71", x"FE", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"FA", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"FE", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"26", x"61", x"16", x"D0", x"18", x"71", x"FE", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"FA", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"FE", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"1C", x"61", x"16", x"D0", x"18", x"70", x"02", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"06", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"02", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"12", x"61", x"16", x"D0", x"18", x"70", x"02", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"06", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"70", x"02", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"A4", x"7A", x"80", x"D0", x"80", x"04", x"80", x"04", x"80", x"04", x"F0", x"1E", 
        x"60", x"12", x"61", x"0C", x"D0", x"18", x"71", x"02", x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"06", 
        x"D0", x"18", x"23", x"EA", x"D0", x"18", x"71", x"02", x"D0", x"18", x"23", x"EA", x"7D", x"01", x"4D", x"07", 
        x"6D", x"00", x"23", x"EA", x"12", x"64", x"6F", x"14", x"FF", x"15", x"FF", x"07", x"3F", x"00", x"13", x"EA", 
        x"6F", x"03", x"FF", x"15", x"00", x"EE", x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", 
        x"FF", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"FF", x"80", x"80", x"80", x"80", x"80", 
        x"80", x"80", x"80", x"80", x"FF", x"00", x"00", x"FF", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", 
        x"20", x"FF", x"38", x"30", x"33", x"33", x"30", x"38", x"3E", x"3C", x"39", x"FF", x"20", x"20", x"20", x"20", 
        x"20", x"20", x"20", x"20", x"20", x"FF", x"00", x"00", x"FF", x"08", x"08", x"08", x"08", x"08", x"08", x"08", 
        x"08", x"08", x"FF", x"38", x"18", x"98", x"98", x"18", x"18", x"38", x"78", x"F8", x"FF", x"08", x"08", x"08", 
        x"08", x"08", x"08", x"08", x"08", x"08", x"FF", x"00", x"00", x"FE", x"02", x"02", x"02", x"02", x"02", x"02", 
        x"02", x"02", x"02", x"FE", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"FE", x"02", x"02", 
        x"02", x"02", x"02", x"02", x"02", x"02", x"02", x"FE", x"00", x"00", x"7C", x"FE", x"C6", x"C6", x"C6", x"FE", 
        x"7C", x"00", x"7C", x"FE", x"C6", x"C0", x"C6", x"FE", x"7C", x"00", x"FE", x"FE", x"38", x"38", x"38", x"38", 
        x"38", x"00", x"7C", x"FE", x"C6", x"C6", x"C6", x"FE", x"7C", x"00", x"FE", x"FE", x"0C", x"0C", x"CC", x"FC", 
        x"78", x"00", x"7C", x"FE", x"C6", x"FE", x"FE", x"C6", x"C6", x"00", x"C6", x"EE", x"FE", x"FE", x"FE", x"D6", 
        x"C6", x"00"
    );

end package;

package body octojam9title is
end octojam9title;