library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package flags is

    type t_ROM is array (0 to 1017 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"12", x"A0", x"60", x"00", x"E0", x"A1", x"12", x"04", x"70", x"01", x"40", x"10", x"00", x"EE", x"12", x"04", 
        x"FC", x"65", x"22", x"76", x"41", x"00", x"00", x"EE", x"80", x"10", x"22", x"76", x"42", x"00", x"00", x"EE", 
        x"80", x"20", x"22", x"76", x"43", x"00", x"00", x"EE", x"80", x"30", x"22", x"76", x"44", x"00", x"00", x"EE", 
        x"80", x"40", x"22", x"76", x"45", x"00", x"00", x"EE", x"80", x"50", x"22", x"76", x"46", x"00", x"00", x"EE", 
        x"80", x"60", x"22", x"76", x"47", x"00", x"00", x"EE", x"80", x"70", x"22", x"76", x"48", x"00", x"00", x"EE", 
        x"80", x"80", x"22", x"76", x"49", x"00", x"00", x"EE", x"80", x"90", x"22", x"76", x"4A", x"00", x"00", x"EE", 
        x"80", x"A0", x"22", x"76", x"4B", x"00", x"00", x"EE", x"80", x"B0", x"22", x"76", x"4C", x"00", x"00", x"EE", 
        x"80", x"C0", x"22", x"76", x"00", x"EE", x"A5", x"3F", x"F0", x"1E", x"DD", x"E4", x"7D", x"04", x"00", x"EE", 
        x"A5", x"43", x"8E", x"D0", x"8E", x"EE", x"8E", x"EE", x"FE", x"1E", x"DA", x"B4", x"7A", x"05", x"00", x"EE", 
        x"A5", x"40", x"92", x"C0", x"A5", x"3D", x"7B", x"01", x"DA", x"B3", x"7A", x"04", x"7B", x"FF", x"00", x"EE", 
        x"00", x"E0", x"6A", x"32", x"6B", x"1B", x"A5", x"F1", x"DA", x"B4", x"6A", x"3A", x"A5", x"F5", x"DA", x"B4", 
        x"6D", x"00", x"6E", x"00", x"A5", x"DF", x"22", x"10", x"6A", x"16", x"6B", x"00", x"61", x"0F", x"6D", x"01", 
        x"22", x"80", x"63", x"0F", x"6F", x"14", x"83", x"F1", x"6F", x"00", x"62", x"32", x"82", x"11", x"8E", x"F0", 
        x"6C", x"3F", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", x"6C", x"1F", x"22", x"90", 
        x"7A", x"05", x"6D", x"02", x"22", x"80", x"63", x"0F", x"6F", x"14", x"83", x"F2", x"6F", x"00", x"62", x"32", 
        x"82", x"12", x"8E", x"F0", x"6C", x"02", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", 
        x"6C", x"04", x"22", x"90", x"7B", x"05", x"6A", x"00", x"6D", x"03", x"22", x"80", x"63", x"0F", x"6F", x"14", 
        x"83", x"F3", x"6F", x"00", x"62", x"32", x"82", x"13", x"8E", x"F0", x"6C", x"3D", x"22", x"90", x"82", x"E0", 
        x"6C", x"00", x"22", x"90", x"82", x"30", x"6C", x"1B", x"22", x"90", x"7A", x"05", x"6D", x"04", x"22", x"80", 
        x"6F", x"14", x"8F", x"14", x"84", x"F0", x"63", x"0F", x"6F", x"14", x"83", x"F4", x"6F", x"AA", x"62", x"32", 
        x"82", x"14", x"8E", x"F0", x"6C", x"41", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", 
        x"6C", x"23", x"22", x"90", x"82", x"40", x"6C", x"00", x"22", x"90", x"7A", x"01", x"6D", x"05", x"22", x"80", 
        x"6F", x"14", x"8F", x"15", x"84", x"F0", x"63", x"14", x"6F", x"0F", x"83", x"F5", x"6F", x"AA", x"62", x"32", 
        x"82", x"15", x"8E", x"F0", x"6C", x"23", x"22", x"90", x"82", x"E0", x"6C", x"01", x"22", x"90", x"82", x"30", 
        x"6C", x"05", x"22", x"90", x"82", x"40", x"6C", x"01", x"22", x"90", x"7B", x"05", x"6A", x"00", x"6D", x"06", 
        x"22", x"80", x"6F", x"3C", x"8F", x"F6", x"83", x"F0", x"6F", x"AA", x"62", x"3C", x"82", x"26", x"8E", x"F0", 
        x"6C", x"1E", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", x"6C", x"00", x"22", x"90", 
        x"7A", x"05", x"6D", x"07", x"22", x"80", x"6F", x"0A", x"8F", x"17", x"84", x"F0", x"63", x"0F", x"6F", x"14", 
        x"83", x"F7", x"6F", x"AA", x"62", x"0F", x"61", x"32", x"82", x"17", x"8E", x"F0", x"6C", x"23", x"22", x"90", 
        x"82", x"E0", x"6C", x"01", x"22", x"90", x"82", x"30", x"6C", x"05", x"22", x"90", x"82", x"40", x"6C", x"01", 
        x"22", x"90", x"7A", x"01", x"6D", x"0E", x"22", x"80", x"6F", x"32", x"8F", x"FE", x"83", x"F0", x"6F", x"AA", 
        x"62", x"32", x"82", x"2E", x"8E", x"F0", x"6C", x"64", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", 
        x"82", x"30", x"6C", x"00", x"22", x"90", x"6D", x"00", x"6E", x"10", x"A5", x"E5", x"22", x"10", x"6A", x"16", 
        x"6B", x"10", x"61", x"64", x"6D", x"04", x"22", x"80", x"6F", x"C8", x"8F", x"14", x"84", x"F0", x"63", x"64", 
        x"6F", x"C8", x"83", x"F4", x"6F", x"AA", x"62", x"C8", x"82", x"14", x"8E", x"F0", x"6C", x"2C", x"22", x"90", 
        x"82", x"E0", x"6C", x"01", x"22", x"90", x"82", x"30", x"6C", x"2C", x"22", x"90", x"82", x"40", x"6C", x"01", 
        x"22", x"90", x"7A", x"01", x"6D", x"05", x"22", x"80", x"6F", x"5F", x"8F", x"15", x"84", x"F0", x"63", x"5F", 
        x"6F", x"64", x"83", x"F5", x"6F", x"AA", x"62", x"5F", x"82", x"15", x"8E", x"F0", x"6C", x"FB", x"22", x"90", 
        x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", x"6C", x"FB", x"22", x"90", x"82", x"40", x"6C", x"00", 
        x"22", x"90", x"7B", x"05", x"6A", x"00", x"6D", x"06", x"22", x"80", x"6F", x"3D", x"8F", x"F6", x"83", x"F0", 
        x"6F", x"AA", x"62", x"3D", x"82", x"26", x"8E", x"F0", x"6C", x"1E", x"22", x"90", x"82", x"E0", x"6C", x"01", 
        x"22", x"90", x"82", x"30", x"6C", x"01", x"22", x"90", x"7A", x"05", x"6D", x"07", x"22", x"80", x"6F", x"69", 
        x"8F", x"17", x"84", x"F0", x"63", x"69", x"6F", x"64", x"83", x"F7", x"6F", x"AA", x"62", x"69", x"82", x"17", 
        x"8E", x"F0", x"6C", x"FB", x"22", x"90", x"82", x"E0", x"6C", x"00", x"22", x"90", x"82", x"30", x"6C", x"FB", 
        x"22", x"90", x"82", x"40", x"6C", x"00", x"22", x"90", x"7A", x"01", x"6D", x"0E", x"22", x"80", x"6F", x"BC", 
        x"8F", x"FE", x"83", x"F0", x"6F", x"AA", x"62", x"BC", x"82", x"2E", x"8E", x"F0", x"6C", x"78", x"22", x"90", 
        x"82", x"E0", x"6C", x"01", x"22", x"90", x"82", x"30", x"6C", x"01", x"22", x"90", x"6D", x"00", x"6E", x"1B", 
        x"A5", x"EB", x"22", x"10", x"6A", x"16", x"6B", x"1B", x"6D", x"0F", x"22", x"80", x"7A", x"FF", x"6D", x"0E", 
        x"22", x"80", x"A5", x"2C", x"61", x"10", x"F1", x"1E", x"60", x"AA", x"F0", x"55", x"A5", x"3C", x"F0", x"65", 
        x"82", x"00", x"6C", x"AA", x"22", x"90", x"A5", x"2C", x"6F", x"10", x"FF", x"1E", x"60", x"55", x"F0", x"55", 
        x"A5", x"3C", x"F0", x"65", x"82", x"00", x"6C", x"55", x"22", x"90", x"15", x"2A", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A0", x"C0", x"80", 
        x"A0", x"40", x"A0", x"E0", x"A0", x"A0", x"E0", x"C0", x"40", x"40", x"E0", x"E0", x"20", x"C0", x"E0", x"E0", 
        x"60", x"20", x"E0", x"A0", x"E0", x"20", x"20", x"E0", x"C0", x"20", x"C0", x"E0", x"80", x"E0", x"E0", x"E0", 
        x"20", x"20", x"20", x"E0", x"E0", x"A0", x"E0", x"E0", x"E0", x"20", x"E0", x"40", x"A0", x"E0", x"A0", x"C0", 
        x"E0", x"A0", x"E0", x"E0", x"80", x"80", x"E0", x"C0", x"A0", x"A0", x"C0", x"E0", x"C0", x"80", x"E0", x"E0", 
        x"80", x"C0", x"80", x"60", x"80", x"A0", x"60", x"A0", x"E0", x"A0", x"A0", x"E0", x"40", x"40", x"E0", x"60", 
        x"20", x"20", x"C0", x"A0", x"C0", x"A0", x"A0", x"80", x"80", x"80", x"E0", x"E0", x"E0", x"A0", x"A0", x"C0", 
        x"A0", x"A0", x"A0", x"E0", x"A0", x"A0", x"E0", x"C0", x"A0", x"C0", x"80", x"40", x"A0", x"E0", x"60", x"C0", 
        x"A0", x"C0", x"A0", x"60", x"C0", x"20", x"C0", x"E0", x"40", x"40", x"40", x"A0", x"A0", x"A0", x"60", x"A0", 
        x"A0", x"A0", x"40", x"A0", x"A0", x"E0", x"E0", x"A0", x"40", x"A0", x"A0", x"A0", x"A0", x"40", x"40", x"E0", 
        x"60", x"80", x"E0", x"00", x"00", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"40", x"48", 
        x"2C", x"68", x"68", x"8C", x"00", x"34", x"2C", x"70", x"70", x"8C", x"00", x"64", x"78", x"48", x"3C", x"70", 
        x"00", x"0A", x"AE", x"A2", x"42", x"38", x"28", x"28", x"B8"
    );

end package;

package body flags is
end flags;