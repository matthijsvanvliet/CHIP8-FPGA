library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package bc_test is

    type t_ROM is array (0 to 470 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"00", x"E0", x"63", x"00", x"64", x"01", x"65", x"EE", x"35", x"EE", x"13", x"10", x"63", x"00", x"64", x"02", 
        x"65", x"EE", x"66", x"EE", x"55", x"60", x"13", x"10", x"63", x"00", x"64", x"03", x"65", x"EE", x"45", x"FD", 
        x"13", x"10", x"63", x"00", x"64", x"04", x"65", x"EE", x"75", x"01", x"35", x"EF", x"13", x"10", x"63", x"00", 
        x"64", x"05", x"6F", x"01", x"65", x"EE", x"66", x"EF", x"85", x"65", x"3F", x"00", x"13", x"10", x"63", x"00", 
        x"64", x"06", x"6F", x"00", x"65", x"EF", x"66", x"EE", x"85", x"65", x"3F", x"01", x"13", x"10", x"6F", x"00", 
        x"63", x"00", x"64", x"07", x"65", x"EE", x"66", x"EF", x"85", x"67", x"3F", x"01", x"13", x"10", x"63", x"00", 
        x"64", x"08", x"6F", x"01", x"65", x"EF", x"66", x"EE", x"85", x"67", x"3F", x"00", x"13", x"10", x"63", x"00", 
        x"64", x"09", x"65", x"F0", x"66", x"0F", x"85", x"61", x"35", x"FF", x"13", x"10", x"63", x"01", x"64", x"00", 
        x"65", x"F0", x"66", x"0F", x"85", x"62", x"35", x"00", x"13", x"10", x"63", x"01", x"64", x"01", x"65", x"F0", 
        x"66", x"0F", x"85", x"63", x"35", x"FF", x"13", x"10", x"6F", x"00", x"63", x"01", x"64", x"02", x"65", x"81", 
        x"85", x"0E", x"3F", x"01", x"13", x"10", x"63", x"01", x"64", x"03", x"6F", x"01", x"65", x"47", x"85", x"0E", 
        x"3F", x"00", x"13", x"10", x"63", x"01", x"64", x"04", x"6F", x"00", x"65", x"01", x"85", x"06", x"3F", x"01", 
        x"13", x"10", x"63", x"01", x"64", x"05", x"6F", x"01", x"65", x"02", x"85", x"06", x"3F", x"00", x"13", x"10", 
        x"63", x"01", x"64", x"06", x"60", x"15", x"61", x"78", x"A3", x"D0", x"F1", x"55", x"F1", x"65", x"30", x"15", 
        x"13", x"10", x"31", x"78", x"13", x"10", x"63", x"01", x"64", x"07", x"60", x"8A", x"A3", x"D0", x"F0", x"33", 
        x"A3", x"D0", x"F0", x"65", x"30", x"01", x"13", x"10", x"60", x"01", x"F0", x"1E", x"F0", x"65", x"30", x"03", 
        x"13", x"10", x"60", x"01", x"F0", x"1E", x"F0", x"65", x"30", x"08", x"13", x"10", x"13", x"32", x"13", x"0E", 
        x"A3", x"2A", x"60", x"13", x"61", x"09", x"D0", x"18", x"F3", x"29", x"60", x"22", x"61", x"0B", x"D0", x"15", 
        x"F4", x"29", x"60", x"28", x"61", x"0B", x"D0", x"15", x"13", x"0E", x"FF", x"F0", x"F0", x"FF", x"F0", x"F0", 
        x"F0", x"FF", x"A3", x"58", x"60", x"15", x"61", x"0B", x"63", x"08", x"D0", x"18", x"70", x"08", x"F3", x"1E", 
        x"30", x"2D", x"13", x"3A", x"A3", x"70", x"60", x"02", x"61", x"18", x"63", x"08", x"D0", x"18", x"70", x"05", 
        x"F3", x"1E", x"30", x"3E", x"13", x"4C", x"13", x"0E", x"F0", x"88", x"88", x"F0", x"88", x"88", x"88", x"F0", 
        x"78", x"84", x"84", x"84", x"84", x"84", x"84", x"78", x"84", x"C4", x"A4", x"94", x"8C", x"84", x"84", x"84", 
        x"C0", x"A0", x"A0", x"C0", x"A0", x"A0", x"C0", x"00", x"00", x"00", x"A0", x"A0", x"E0", x"20", x"20", x"E0", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"C0", x"A0", x"A0", x"C0", x"A0", x"A0", x"C0", x"00", 
        x"00", x"00", x"60", x"A0", x"C0", x"80", x"60", x"00", x"00", x"00", x"60", x"80", x"40", x"20", x"C0", x"00", 
        x"80", x"80", x"C0", x"80", x"80", x"80", x"60", x"00", x"E0", x"80", x"80", x"80", x"80", x"80", x"E0", x"00", 
        x"00", x"00", x"40", x"A0", x"A0", x"A0", x"40", x"00", x"20", x"20", x"20", x"60", x"A0", x"A0", x"60", x"00", 
        x"00", x"00", x"60", x"A0", x"C0", x"80", x"60", x"00", x"00", x"00", x"00", x"60", x"40", x"40", x"50", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00"
    );

end package;

package body bc_test is
end bc_test;