library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package keypad_test is

    type t_ROM is array (0 to 913 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"13", x"0C", x"60", x"00", x"E0", x"A1", x"12", x"04", x"70", x"01", x"40", x"10", x"00", x"EE", x"12", x"04", 
        x"65", x"00", x"A2", x"22", x"F1", x"55", x"A2", x"82", x"F1", x"55", x"12", x"22", x"43", x"01", x"D0", x"12", 
        x"22", x"02", x"00", x"00", x"F5", x"1E", x"F5", x"1E", x"F5", x"1E", x"F5", x"1E", x"F1", x"65", x"63", x"00", 
        x"F3", x"15", x"F4", x"07", x"34", x"00", x"12", x"44", x"A4", x"23", x"D0", x"12", x"64", x"0A", x"F4", x"15", 
        x"64", x"01", x"83", x"43", x"64", x"0E", x"E4", x"9E", x"12", x"52", x"45", x"00", x"12", x"52", x"75", x"FF", 
        x"12", x"1C", x"64", x"0F", x"E4", x"9E", x"12", x"60", x"95", x"20", x"12", x"60", x"75", x"01", x"12", x"1C", 
        x"86", x"50", x"64", x"0A", x"E4", x"A1", x"12", x"80", x"64", x"00", x"72", x"01", x"74", x"01", x"E4", x"9E", 
        x"12", x"78", x"86", x"40", x"76", x"FF", x"12", x"80", x"54", x"20", x"12", x"6C", x"72", x"FF", x"12", x"32", 
        x"22", x"02", x"00", x"00", x"F6", x"1E", x"F6", x"1E", x"F6", x"1E", x"F6", x"1E", x"64", x"02", x"F4", x"1E", 
        x"F1", x"65", x"64", x"10", x"80", x"41", x"A2", x"9A", x"F1", x"55", x"00", x"00", x"FC", x"65", x"23", x"02", 
        x"41", x"00", x"00", x"EE", x"80", x"10", x"23", x"02", x"42", x"00", x"00", x"EE", x"80", x"20", x"23", x"02", 
        x"43", x"00", x"00", x"EE", x"80", x"30", x"23", x"02", x"44", x"00", x"00", x"EE", x"80", x"40", x"23", x"02", 
        x"45", x"00", x"00", x"EE", x"80", x"50", x"23", x"02", x"46", x"00", x"00", x"EE", x"80", x"60", x"23", x"02", 
        x"47", x"00", x"00", x"EE", x"80", x"70", x"23", x"02", x"48", x"00", x"00", x"EE", x"80", x"80", x"23", x"02", 
        x"49", x"00", x"00", x"EE", x"80", x"90", x"23", x"02", x"4A", x"00", x"00", x"EE", x"80", x"A0", x"23", x"02", 
        x"4B", x"00", x"00", x"EE", x"80", x"B0", x"23", x"02", x"4C", x"00", x"00", x"EE", x"80", x"C0", x"23", x"02", 
        x"00", x"EE", x"A4", x"27", x"F0", x"1E", x"DD", x"E4", x"7D", x"04", x"00", x"EE", x"00", x"E0", x"A1", x"FF", 
        x"F0", x"65", x"40", x"01", x"13", x"54", x"40", x"02", x"13", x"58", x"40", x"03", x"13", x"BE", x"6D", x"0A", 
        x"6E", x"02", x"A4", x"D3", x"22", x"9C", x"6D", x"08", x"6E", x"0A", x"A4", x"DF", x"22", x"9C", x"6D", x"08", 
        x"6E", x"0F", x"A4", x"EB", x"22", x"9C", x"6D", x"08", x"6E", x"14", x"A4", x"F5", x"22", x"9C", x"6A", x"32", 
        x"6B", x"1B", x"A5", x"89", x"DA", x"B4", x"6A", x"3A", x"A5", x"8D", x"DA", x"B4", x"60", x"A4", x"61", x"C7", 
        x"62", x"02", x"12", x"10", x"61", x"9E", x"13", x"5A", x"61", x"A1", x"60", x"EE", x"A3", x"9E", x"F1", x"55", 
        x"00", x"E0", x"A5", x"33", x"FF", x"65", x"A4", x"12", x"FF", x"55", x"6D", x"12", x"6E", x"03", x"A5", x"43", 
        x"22", x"9C", x"6D", x"12", x"6E", x"0A", x"A5", x"4B", x"22", x"9C", x"6D", x"12", x"6E", x"11", x"A5", x"53", 
        x"22", x"9C", x"6D", x"12", x"6E", x"18", x"A5", x"5B", x"22", x"9C", x"6E", x"00", x"23", x"96", x"7E", x"01", 
        x"4E", x"10", x"6E", x"00", x"13", x"8C", x"A4", x"12", x"FE", x"1E", x"F0", x"65", x"62", x"01", x"EE", x"A1", 
        x"62", x"00", x"90", x"20", x"13", x"BC", x"80", x"E0", x"80", x"0E", x"A5", x"63", x"F0", x"1E", x"F1", x"65", 
        x"A5", x"83", x"D0", x"16", x"A4", x"12", x"FE", x"1E", x"80", x"20", x"F0", x"55", x"00", x"EE", x"00", x"E0", 
        x"6D", x"06", x"6E", x"0D", x"A5", x"03", x"22", x"9C", x"60", x"03", x"F0", x"15", x"F0", x"0A", x"F1", x"07", 
        x"31", x"00", x"13", x"F2", x"E0", x"A1", x"13", x"F8", x"00", x"E0", x"A4", x"25", x"60", x"1E", x"61", x"09", 
        x"D0", x"13", x"6D", x"10", x"6E", x"11", x"A5", x"11", x"22", x"9C", x"22", x"02", x"F0", x"0A", x"22", x"02", 
        x"13", x"0C", x"6D", x"0A", x"A5", x"1A", x"13", x"FC", x"6D", x"08", x"A5", x"26", x"00", x"E0", x"6E", x"11", 
        x"22", x"9C", x"A4", x"28", x"60", x"1E", x"61", x"09", x"D0", x"13", x"22", x"02", x"F0", x"0A", x"22", x"02", 
        x"13", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"C0", x"C0", x"A0", x"C0", x"80", x"A0", x"40", x"A0", x"E0", x"A0", x"A0", x"E0", x"C0", 
        x"40", x"40", x"E0", x"E0", x"20", x"C0", x"E0", x"E0", x"60", x"20", x"E0", x"A0", x"E0", x"20", x"20", x"E0", 
        x"C0", x"20", x"C0", x"E0", x"80", x"E0", x"E0", x"E0", x"20", x"20", x"20", x"E0", x"E0", x"A0", x"E0", x"E0", 
        x"E0", x"20", x"E0", x"40", x"A0", x"E0", x"A0", x"C0", x"E0", x"A0", x"E0", x"E0", x"80", x"80", x"E0", x"C0", 
        x"A0", x"A0", x"C0", x"E0", x"C0", x"80", x"E0", x"E0", x"80", x"C0", x"80", x"60", x"80", x"A0", x"60", x"A0", 
        x"E0", x"A0", x"A0", x"E0", x"40", x"40", x"E0", x"60", x"20", x"20", x"C0", x"A0", x"C0", x"A0", x"A0", x"80", 
        x"80", x"80", x"E0", x"E0", x"E0", x"A0", x"A0", x"C0", x"A0", x"A0", x"A0", x"E0", x"A0", x"A0", x"E0", x"C0", 
        x"A0", x"C0", x"80", x"40", x"A0", x"E0", x"60", x"C0", x"A0", x"C0", x"A0", x"60", x"C0", x"20", x"C0", x"E0", 
        x"40", x"40", x"40", x"A0", x"A0", x"A0", x"60", x"A0", x"A0", x"A0", x"40", x"A0", x"A0", x"E0", x"E0", x"A0", 
        x"40", x"A0", x"A0", x"A0", x"A0", x"40", x"40", x"E0", x"60", x"80", x"E0", x"00", x"00", x"00", x"00", x"00", 
        x"E0", x"00", x"00", x"00", x"00", x"00", x"40", x"04", x"0B", x"03", x"54", x"04", x"10", x"03", x"58", x"04", 
        x"15", x"03", x"BE", x"68", x"4C", x"34", x"54", x"94", x"64", x"68", x"34", x"64", x"38", x"3C", x"00", x"08", 
        x"94", x"3C", x"88", x"28", x"3C", x"94", x"38", x"64", x"84", x"60", x"00", x"0C", x"94", x"3C", x"88", x"2C", 
        x"08", x"94", x"7C", x"68", x"00", x"10", x"94", x"40", x"88", x"04", x"2C", x"94", x"44", x"3C", x"78", x"54", 
        x"3C", x"8C", x"00", x"68", x"70", x"3C", x"74", x"74", x"94", x"2C", x"60", x"8C", x"94", x"54", x"3C", x"8C", 
        x"00", x"2C", x"58", x"58", x"94", x"44", x"64", x"64", x"38", x"00", x"60", x"64", x"78", x"94", x"48", x"2C", 
        x"58", x"78", x"4C", x"60", x"44", x"00", x"60", x"64", x"78", x"94", x"70", x"3C", x"58", x"3C", x"2C", x"74", 
        x"3C", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"08", x"94", x"0C", x"94", x"10", x"94", x"34", x"00", x"14", x"94", x"18", x"94", x"1C", 
        x"94", x"38", x"00", x"20", x"94", x"24", x"94", x"28", x"94", x"3C", x"00", x"2C", x"94", x"04", x"94", x"30", 
        x"94", x"40", x"00", x"18", x"17", x"10", x"02", x"18", x"02", x"20", x"02", x"10", x"09", x"18", x"09", x"20", 
        x"09", x"10", x"10", x"18", x"10", x"20", x"10", x"10", x"17", x"20", x"17", x"28", x"02", x"28", x"09", x"28", 
        x"10", x"28", x"17", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"0A", x"AE", x"A2", x"42", x"38", x"28", x"28", 
        x"B8"
    );

end package;

package body keypad_test is
end keypad_test;