library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package spaceinvaders is

    type t_ROM is array (0 to 1301 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"12", x"25", x"53", x"50", x"41", x"43", x"45", x"20", x"49", x"4E", x"56", x"41", x"44", x"45", x"52", x"53", 
        x"20", x"30", x"2E", x"39", x"31", x"20", x"42", x"79", x"20", x"44", x"61", x"76", x"69", x"64", x"20", x"57", 
        x"49", x"4E", x"54", x"45", x"52", x"60", x"00", x"61", x"00", x"62", x"08", x"A3", x"DD", x"D0", x"18", x"71", 
        x"08", x"F2", x"1E", x"31", x"20", x"12", x"2D", x"70", x"08", x"61", x"00", x"30", x"40", x"12", x"2D", x"69", 
        x"05", x"6C", x"15", x"6E", x"00", x"23", x"91", x"60", x"0A", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", 
        x"4B", x"23", x"91", x"7E", x"01", x"12", x"45", x"66", x"00", x"68", x"1C", x"69", x"00", x"6A", x"04", x"6B", 
        x"0A", x"6C", x"04", x"6D", x"3C", x"6E", x"0F", x"00", x"E0", x"23", x"75", x"23", x"51", x"FD", x"15", x"60", 
        x"04", x"E0", x"9E", x"12", x"7D", x"23", x"75", x"38", x"00", x"78", x"FF", x"23", x"75", x"60", x"06", x"E0", 
        x"9E", x"12", x"8B", x"23", x"75", x"38", x"39", x"78", x"01", x"23", x"75", x"36", x"00", x"12", x"9F", x"60", 
        x"05", x"E0", x"9E", x"12", x"E9", x"66", x"01", x"65", x"1B", x"84", x"80", x"A3", x"D9", x"D4", x"51", x"A3", 
        x"D9", x"D4", x"51", x"75", x"FF", x"35", x"FF", x"12", x"AD", x"66", x"00", x"12", x"E9", x"D4", x"51", x"3F", 
        x"01", x"12", x"E9", x"D4", x"51", x"66", x"00", x"83", x"40", x"73", x"03", x"83", x"B5", x"62", x"F8", x"83", 
        x"22", x"62", x"08", x"33", x"00", x"12", x"C9", x"23", x"7D", x"82", x"06", x"43", x"08", x"12", x"D3", x"33", 
        x"10", x"12", x"D5", x"23", x"7D", x"82", x"06", x"33", x"18", x"12", x"DD", x"23", x"7D", x"82", x"06", x"43", 
        x"20", x"12", x"E7", x"33", x"28", x"12", x"E9", x"23", x"7D", x"3E", x"00", x"13", x"07", x"79", x"06", x"49", 
        x"18", x"69", x"00", x"6A", x"04", x"6B", x"0A", x"6C", x"04", x"7D", x"F4", x"6E", x"0F", x"00", x"E0", x"23", 
        x"51", x"23", x"75", x"FD", x"15", x"12", x"6F", x"F7", x"07", x"37", x"00", x"12", x"6F", x"FD", x"15", x"23", 
        x"51", x"8B", x"A4", x"3B", x"12", x"13", x"1B", x"7C", x"02", x"6A", x"FC", x"3B", x"02", x"13", x"23", x"7C", 
        x"02", x"6A", x"04", x"23", x"51", x"3C", x"18", x"12", x"6F", x"00", x"E0", x"A4", x"DD", x"60", x"14", x"61", 
        x"08", x"62", x"0F", x"D0", x"1F", x"70", x"08", x"F2", x"1E", x"30", x"2C", x"13", x"33", x"60", x"FF", x"F0", 
        x"15", x"F0", x"07", x"30", x"00", x"13", x"41", x"F0", x"0A", x"00", x"E0", x"A7", x"06", x"FE", x"65", x"12", 
        x"25", x"A3", x"C1", x"F9", x"1E", x"61", x"08", x"23", x"69", x"81", x"06", x"23", x"69", x"81", x"06", x"23", 
        x"69", x"81", x"06", x"23", x"69", x"7B", x"D0", x"00", x"EE", x"80", x"E0", x"80", x"12", x"30", x"00", x"DB", 
        x"C6", x"7B", x"0C", x"00", x"EE", x"A3", x"D9", x"60", x"1C", x"D8", x"04", x"00", x"EE", x"23", x"51", x"8E", 
        x"23", x"23", x"51", x"60", x"05", x"F0", x"18", x"F0", x"15", x"F0", x"07", x"30", x"00", x"13", x"89", x"00", 
        x"EE", x"6A", x"00", x"8D", x"E0", x"6B", x"04", x"E9", x"A1", x"12", x"57", x"A6", x"0C", x"FD", x"1E", x"F0", 
        x"65", x"30", x"FF", x"13", x"AF", x"6A", x"00", x"6B", x"04", x"6D", x"01", x"6E", x"01", x"13", x"97", x"A5", 
        x"0A", x"F0", x"1E", x"DB", x"C6", x"7B", x"08", x"7D", x"01", x"7A", x"01", x"3A", x"07", x"13", x"97", x"00", 
        x"EE", x"3C", x"7E", x"FF", x"FF", x"99", x"99", x"7E", x"FF", x"FF", x"24", x"24", x"E7", x"7E", x"FF", x"3C", 
        x"3C", x"7E", x"DB", x"81", x"42", x"3C", x"7E", x"FF", x"DB", x"10", x"38", x"7C", x"FE", x"00", x"00", x"7F", 
        x"00", x"3F", x"00", x"7F", x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"00", x"00", 
        x"3F", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"3F", x"08", x"08", x"FF", x"00", x"00", x"FE", 
        x"00", x"FC", x"00", x"FE", x"00", x"00", x"00", x"7E", x"42", x"42", x"62", x"62", x"62", x"62", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"7D", x"00", 
        x"41", x"7D", x"05", x"7D", x"7D", x"00", x"00", x"C2", x"C2", x"C6", x"44", x"6C", x"28", x"38", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"F7", x"10", 
        x"14", x"F7", x"F7", x"04", x"04", x"00", x"00", x"7C", x"44", x"FE", x"C2", x"C2", x"C2", x"C2", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"EF", x"20", 
        x"28", x"E8", x"E8", x"2F", x"2F", x"00", x"00", x"F9", x"85", x"C5", x"C5", x"C5", x"C5", x"F9", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"BE", x"00", 
        x"20", x"30", x"20", x"BE", x"BE", x"00", x"00", x"F7", x"04", x"E7", x"85", x"85", x"84", x"F4", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"7F", 
        x"00", x"3F", x"00", x"7F", x"00", x"00", x"00", x"EF", x"28", x"EF", x"00", x"E0", x"60", x"6F", x"00", x"00", 
        x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FE", 
        x"00", x"FC", x"00", x"FE", x"00", x"00", x"00", x"C0", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", 
        x"FC", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"04", x"FC", x"10", x"10", x"FF", x"F9", x"81", x"B9", 
        x"8B", x"9A", x"9A", x"FA", x"00", x"FA", x"8A", x"9A", x"9A", x"9B", x"99", x"F8", x"E6", x"25", x"25", x"F4", 
        x"34", x"34", x"34", x"00", x"17", x"14", x"34", x"37", x"36", x"26", x"C7", x"DF", x"50", x"50", x"5C", x"D8", 
        x"D8", x"DF", x"00", x"DF", x"11", x"1F", x"12", x"1B", x"19", x"D9", x"7C", x"44", x"FE", x"86", x"86", x"86", 
        x"FC", x"84", x"FE", x"82", x"82", x"FE", x"FE", x"80", x"C0", x"C0", x"C0", x"FE", x"FC", x"82", x"C2", x"C2", 
        x"C2", x"FC", x"FE", x"80", x"F8", x"C0", x"C0", x"FE", x"FE", x"80", x"F0", x"C0", x"C0", x"C0", x"FE", x"80", 
        x"BE", x"86", x"86", x"FE", x"86", x"86", x"FE", x"86", x"86", x"86", x"10", x"10", x"10", x"10", x"10", x"10", 
        x"18", x"18", x"18", x"48", x"48", x"78", x"9C", x"90", x"B0", x"C0", x"B0", x"9C", x"80", x"80", x"C0", x"C0", 
        x"C0", x"FE", x"EE", x"92", x"92", x"86", x"86", x"86", x"FE", x"82", x"86", x"86", x"86", x"86", x"7C", x"82", 
        x"86", x"86", x"86", x"7C", x"FE", x"82", x"FE", x"C0", x"C0", x"C0", x"7C", x"82", x"C2", x"CA", x"C4", x"7A", 
        x"FE", x"86", x"FE", x"90", x"9C", x"84", x"FE", x"C0", x"FE", x"02", x"02", x"FE", x"FE", x"10", x"30", x"30", 
        x"30", x"30", x"82", x"82", x"C2", x"C2", x"C2", x"FE", x"82", x"82", x"82", x"EE", x"38", x"10", x"86", x"86", 
        x"96", x"92", x"92", x"EE", x"82", x"44", x"38", x"38", x"44", x"82", x"82", x"82", x"FE", x"30", x"30", x"30", 
        x"FE", x"02", x"1E", x"F0", x"80", x"FE", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"00", x"00", x"60", 
        x"60", x"C0", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"18", x"00", x"18", x"7C", x"C6", 
        x"0C", x"18", x"00", x"18", x"00", x"00", x"FE", x"FE", x"00", x"00", x"FE", x"82", x"86", x"86", x"86", x"FE", 
        x"08", x"08", x"08", x"18", x"18", x"18", x"FE", x"02", x"FE", x"C0", x"C0", x"FE", x"FE", x"02", x"1E", x"06", 
        x"06", x"FE", x"84", x"C4", x"C4", x"FE", x"04", x"04", x"FE", x"80", x"FE", x"06", x"06", x"FE", x"C0", x"C0", 
        x"C0", x"FE", x"82", x"FE", x"FE", x"02", x"02", x"06", x"06", x"06", x"7C", x"44", x"FE", x"86", x"86", x"FE", 
        x"FE", x"82", x"FE", x"06", x"06", x"06", x"44", x"FE", x"44", x"44", x"FE", x"44", x"A8", x"A8", x"A8", x"A8", 
        x"A8", x"A8", x"A8", x"6C", x"5A", x"00", x"0C", x"18", x"A8", x"30", x"4E", x"7E", x"00", x"12", x"18", x"66", 
        x"6C", x"A8", x"5A", x"66", x"54", x"24", x"66", x"00", x"48", x"48", x"18", x"12", x"A8", x"06", x"90", x"A8", 
        x"12", x"00", x"7E", x"30", x"12", x"A8", x"84", x"30", x"4E", x"72", x"18", x"66", x"A8", x"A8", x"A8", x"A8", 
        x"A8", x"A8", x"90", x"54", x"78", x"A8", x"48", x"78", x"6C", x"72", x"A8", x"12", x"18", x"6C", x"72", x"66", 
        x"54", x"90", x"A8", x"72", x"2A", x"18", x"A8", x"30", x"4E", x"7E", x"00", x"12", x"18", x"66", x"6C", x"A8", 
        x"72", x"54", x"A8", x"5A", x"66", x"18", x"7E", x"18", x"4E", x"72", x"A8", x"72", x"2A", x"18", x"30", x"66", 
        x"A8", x"30", x"4E", x"7E", x"00", x"6C", x"30", x"54", x"4E", x"9C", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
        x"A8", x"48", x"54", x"7E", x"18", x"A8", x"90", x"54", x"78", x"66", x"A8", x"6C", x"2A", x"30", x"5A", x"A8", 
        x"84", x"30", x"72", x"2A", x"A8", x"D8", x"A8", x"00", x"4E", x"12", x"A8", x"E4", x"A2", x"A8", x"00", x"4E", 
        x"12", x"A8", x"6C", x"2A", x"54", x"54", x"72", x"A8", x"84", x"30", x"72", x"2A", x"A8", x"DE", x"9C", x"A8", 
        x"72", x"2A", x"18", x"A8", x"0C", x"54", x"48", x"5A", x"78", x"72", x"18", x"66", x"A8", x"66", x"18", x"5A", 
        x"54", x"66", x"72", x"6C", x"A8", x"72", x"2A", x"00", x"72", x"A8", x"72", x"2A", x"18", x"A8", x"30", x"4E", 
        x"7E", x"00", x"12", x"18", x"66", x"6C", x"A8", x"00", x"66", x"18", x"A8", x"30", x"4E", x"0C", x"66", x"18", 
        x"00", x"6C", x"30", x"4E", x"24", x"A8", x"72", x"2A", x"18", x"30", x"66", x"A8", x"1E", x"54", x"66", x"0C", 
        x"18", x"9C", x"A8", x"24", x"54", x"54", x"12", x"A8", x"42", x"78", x"0C", x"3C", x"A8", x"AE", x"A8", x"A8", 
        x"A8", x"A8", x"A8", x"A8", x"A8", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00"
    );

end package;

package body spaceinvaders is
end spaceinvaders;