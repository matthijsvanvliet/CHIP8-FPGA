library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package sctest is

    type t_ROM is array (0 to 672 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"12", x"12", x"20", x"54", x"72", x"6F", x"6E", x"69", x"78", x"20", x"28", x"63", x"29", x"20", x"32", x"30", 
        x"31", x"30", x"00", x"E0", x"3F", x"00", x"13", x"E2", x"3E", x"00", x"13", x"E2", x"3D", x"00", x"13", x"E2", 
        x"3C", x"00", x"13", x"E2", x"3B", x"00", x"13", x"E2", x"3A", x"00", x"13", x"E2", x"39", x"00", x"13", x"E2", 
        x"38", x"00", x"13", x"E2", x"37", x"00", x"13", x"E2", x"36", x"00", x"13", x"E2", x"35", x"00", x"13", x"E2", 
        x"34", x"00", x"13", x"E2", x"33", x"00", x"13", x"E2", x"32", x"00", x"13", x"E2", x"31", x"00", x"13", x"E2", 
        x"30", x"00", x"13", x"E2", x"60", x"00", x"61", x"01", x"62", x"02", x"63", x"03", x"64", x"04", x"65", x"05", 
        x"66", x"06", x"67", x"07", x"68", x"08", x"69", x"09", x"6A", x"0A", x"6B", x"0B", x"6C", x"0C", x"6D", x"0D", 
        x"6E", x"0E", x"6F", x"0F", x"A4", x"78", x"FF", x"65", x"3F", x"00", x"13", x"F8", x"3E", x"00", x"13", x"F8", 
        x"3D", x"00", x"13", x"F8", x"3C", x"00", x"13", x"F8", x"3B", x"00", x"13", x"F8", x"3A", x"00", x"13", x"F8", 
        x"39", x"00", x"13", x"F8", x"38", x"00", x"13", x"F8", x"37", x"00", x"13", x"F8", x"36", x"00", x"13", x"F8", 
        x"35", x"00", x"13", x"F8", x"34", x"00", x"13", x"F8", x"33", x"00", x"13", x"F8", x"32", x"00", x"13", x"F8", 
        x"31", x"00", x"13", x"F8", x"30", x"00", x"13", x"F8", x"60", x"00", x"F0", x"29", x"F0", x"65", x"40", x"00", 
        x"14", x"02", x"A4", x"52", x"6E", x"7B", x"FE", x"33", x"F2", x"65", x"30", x"01", x"13", x"C6", x"31", x"02", 
        x"13", x"C6", x"32", x"03", x"13", x"C6", x"6E", x"02", x"6F", x"00", x"60", x"FE", x"61", x"01", x"80", x"14", 
        x"3F", x"00", x"14", x"0C", x"6E", x"03", x"30", x"FF", x"14", x"0C", x"6E", x"04", x"80", x"14", x"3F", x"01", 
        x"14", x"0C", x"6E", x"05", x"30", x"00", x"14", x"0C", x"60", x"01", x"6E", x"06", x"6F", x"00", x"80", x"15", 
        x"3F", x"01", x"14", x"0C", x"6E", x"07", x"30", x"00", x"14", x"0C", x"6E", x"08", x"80", x"15", x"3F", x"00", 
        x"14", x"0C", x"6E", x"09", x"30", x"FF", x"14", x"0C", x"60", x"01", x"6E", x"0A", x"6F", x"00", x"80", x"17", 
        x"3F", x"01", x"14", x"0C", x"6E", x"0B", x"30", x"00", x"14", x"0C", x"6E", x"0C", x"60", x"01", x"61", x"00", 
        x"80", x"17", x"3F", x"00", x"14", x"0C", x"6E", x"0D", x"30", x"FF", x"14", x"0C", x"60", x"FF", x"6E", x"0E", 
        x"6F", x"00", x"80", x"06", x"3F", x"01", x"14", x"0C", x"6E", x"0F", x"30", x"7F", x"14", x"0C", x"60", x"40", 
        x"6E", x"10", x"80", x"06", x"3F", x"00", x"14", x"0C", x"6E", x"11", x"30", x"20", x"14", x"0C", x"6E", x"12", 
        x"6F", x"01", x"80", x"0E", x"3F", x"00", x"14", x"0C", x"6E", x"13", x"30", x"40", x"14", x"0C", x"60", x"FA", 
        x"6E", x"14", x"80", x"0E", x"3F", x"01", x"14", x"0C", x"6E", x"15", x"30", x"F4", x"14", x"0C", x"61", x"7B", 
        x"6E", x"16", x"80", x"13", x"30", x"8F", x"14", x"0C", x"A4", x"88", x"F7", x"65", x"F7", x"75", x"A4", x"78", 
        x"F7", x"65", x"F7", x"85", x"6E", x"17", x"37", x"07", x"14", x"0C", x"36", x"06", x"14", x"0C", x"35", x"05", 
        x"14", x"0C", x"34", x"04", x"14", x"0C", x"33", x"03", x"14", x"0C", x"32", x"02", x"14", x"0C", x"31", x"01", 
        x"14", x"0C", x"30", x"00", x"14", x"0C", x"6E", x"18", x"AF", x"FE", x"60", x"02", x"6F", x"00", x"F0", x"1E", 
        x"3F", x"01", x"14", x"0C", x"14", x"90", x"24", x"12", x"70", x"0A", x"62", x"0B", x"F2", x"29", x"D0", x"15", 
        x"70", x"05", x"62", x"0C", x"F2", x"29", x"D0", x"15", x"72", x"01", x"F2", x"29", x"70", x"05", x"D0", x"15", 
        x"14", x"50", x"24", x"12", x"70", x"0A", x"A4", x"64", x"D0", x"15", x"70", x"06", x"A4", x"69", x"D0", x"15", 
        x"70", x"06", x"A4", x"64", x"D0", x"15", x"14", x"50", x"24", x"12", x"70", x"0A", x"A4", x"5A", x"D0", x"15", 
        x"14", x"50", x"24", x"12", x"70", x"0A", x"A4", x"55", x"D0", x"15", x"14", x"50", x"24", x"12", x"24", x"32", 
        x"14", x"50", x"60", x"00", x"61", x"00", x"A4", x"5F", x"D0", x"15", x"70", x"05", x"A4", x"6E", x"D0", x"15", 
        x"70", x"06", x"D0", x"15", x"A4", x"5A", x"70", x"06", x"D0", x"15", x"A4", x"6E", x"70", x"05", x"D0", x"15", 
        x"00", x"EE", x"84", x"00", x"74", x"0A", x"85", x"10", x"A4", x"52", x"FE", x"33", x"F2", x"65", x"F0", x"29", 
        x"D4", x"55", x"74", x"06", x"F1", x"29", x"D4", x"55", x"74", x"06", x"F2", x"29", x"D4", x"55", x"00", x"EE", 
        x"14", x"50", x"00", x"00", x"00", x"10", x"30", x"10", x"10", x"10", x"F0", x"90", x"90", x"90", x"F0", x"F0", 
        x"80", x"F0", x"80", x"F0", x"F8", x"20", x"20", x"20", x"F8", x"88", x"C8", x"A8", x"98", x"88", x"E0", x"90", 
        x"E0", x"90", x"88", x"90", x"A0", x"C0", x"A0", x"90", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"02", x"03", x"04", x"05", x"06", x"07", 
        x"60", x"00", x"61", x"00", x"F0", x"29", x"D0", x"15", x"70", x"05", x"A4", x"73", x"D0", x"15", x"14", x"50"
    );

end package;

package body sctest is
end sctest;