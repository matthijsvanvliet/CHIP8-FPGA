library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package rps is

    type t_ROM is array (0 to 2017 - 1) of std_logic_vector(7 downto 0);
    constant c_ROM : t_ROM := (
        x"17", x"8D", x"3C", x"42", x"A1", x"8B", x"95", x"8B", x"56", x"3C", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"78", x"4C", x"4E", x"42", x"42", x"42", x"42", x"7E", x"00", x"00", x"00", x"00", x"00", x"00", x"C3", x"A5", 
        x"66", x"3C", x"18", x"66", x"C3", x"81", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"9F", x"3F", x"5F", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FC", x"C0", x"FF", x"FF", x"FF", x"7F", x"3F", x"1F", x"0F", x"07", x"FF", x"FF", x"FF", x"FE", 
        x"FC", x"F8", x"F0", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"3F", x"03", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"F9", x"FC", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"03", 
        x"3B", x"C7", x"3F", x"FF", x"7F", x"BF", x"7F", x"00", x"00", x"01", x"1E", x"01", x"00", x"70", x"FD", x"F8", 
        x"88", x"00", x"B0", x"F8", x"00", x"00", x"E0", x"F3", x"73", x"37", x"77", x"E7", x"00", x"00", x"CF", x"EF", 
        x"EE", x"EE", x"CE", x"8F", x"00", x"07", x"8F", x"0F", x"0F", x"1C", x"1D", x"1F", x"FE", x"FD", x"FE", x"00", 
        x"00", x"80", x"78", x"80", x"FF", x"FF", x"FF", x"C0", x"DC", x"E3", x"FC", x"FF", x"FF", x"FF", x"FF", x"1F", 
        x"03", x"FB", x"07", x"FF", x"1F", x"0F", x"01", x"00", x"00", x"FF", x"80", x"7F", x"FC", x"38", x"F8", x"F8", 
        x"E0", x"01", x"00", x"00", x"C3", x"00", x"01", x"03", x"03", x"00", x"00", x"02", x"8F", x"CE", x"EE", x"EE", 
        x"CE", x"8C", x"00", x"40", x"1F", x"1F", x"1D", x"1C", x"1C", x"84", x"00", x"00", x"F8", x"F0", x"80", x"00", 
        x"00", x"FF", x"01", x"FE", x"FF", x"FF", x"FF", x"F8", x"C0", x"DF", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"3F", x"3F", x"9F", x"7F", x"FF", x"FF", x"FF", x"FF", x"E0", x"1C", x"E3", x"FC", 
        x"FF", x"FF", x"FF", x"FF", x"05", x"0A", x"17", x"2F", x"5F", x"BF", x"7F", x"FF", x"A0", x"50", x"E8", x"F4", 
        x"FA", x"FD", x"FE", x"FF", x"07", x"38", x"C7", x"3F", x"FF", x"FF", x"FF", x"FF", x"FC", x"FC", x"F9", x"FE", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"05", x"0B", x"17", x"2F", 
        x"5F", x"BF", x"7F", x"FF", x"E0", x"C0", x"80", x"00", x"00", x"00", x"01", x"00", x"FF", x"FF", x"FF", x"FF", 
        x"FE", x"FC", x"7C", x"FA", x"5F", x"2F", x"17", x"0B", x"05", x"02", x"01", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"F8", x"04", x"06", x"06", x"06", x"06", x"00", x"00", x"1F", x"20", 
        x"20", x"20", x"20", x"20", x"00", x"80", x"40", x"A0", x"D0", x"F0", x"E0", x"C0", x"FD", x"FE", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"07", x"05", x"05", x"05", x"05", x"FF", x"FF", x"FF", x"E0", 
        x"E0", x"E0", x"E0", x"E0", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"FC", x"02", x"06", x"06", x"06", x"06", x"06", x"CE", x"EC", x"1D", x"20", x"20", x"20", x"20", 
        x"20", x"1F", x"0F", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"FF", x"FF", x"FE", x"FC", 
        x"FC", x"FA", x"FD", x"FE", x"05", x"05", x"05", x"05", x"05", x"FD", x"03", x"FF", x"E0", x"E0", x"E0", x"E0", 
        x"E0", x"73", x"36", x"BD", x"FF", x"FF", x"FF", x"FF", x"FF", x"80", x"3F", x"40", x"4A", x"4A", x"02", x"02", 
        x"7A", x"02", x"FC", x"00", x"09", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"40", x"A0", x"D0", x"F0", x"E0", x"C0", x"80", x"00", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"BF", x"BF", x"BF", x"BF", 
        x"BF", x"BF", x"3F", x"7F", x"7F", x"7F", x"40", x"40", x"5E", x"40", x"3F", x"80", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"4F", x"87", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"71", x"75", x"71", 
        x"17", x"FF", x"E9", x"D0", x"FF", x"51", x"17", x"53", x"51", x"FF", x"FF", x"3F", x"FF", x"1F", x"3F", x"DF", 
        x"1F", x"FF", x"FE", x"FD", x"FF", x"11", x"55", x"31", x"57", x"FF", x"DF", x"A7", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F4", x"03", x"01", x"00", x"00", 
        x"00", x"00", x"80", x"00", x"7D", x"3A", x"14", x"08", x"00", x"00", x"BB", x"AA", x"A0", x"40", x"80", x"00", 
        x"00", x"00", x"BB", x"22", x"1F", x"0F", x"06", x"03", x"00", x"00", x"BB", x"12", x"FA", x"F4", x"E8", x"50", 
        x"20", x"00", x"3B", x"A2", x"43", x"81", x"00", x"00", x"00", x"00", x"D5", x"18", x"7F", x"3E", x"1D", x"0A", 
        x"04", x"00", x"DD", x"55", x"E8", x"D0", x"A0", x"40", x"80", x"00", x"01", x"01", x"80", x"80", x"00", x"00", 
        x"E0", x"A0", x"C0", x"A0", x"B1", x"AB", x"00", x"00", x"EE", x"A8", x"EC", x"8E", x"9A", x"BB", x"00", x"00", 
        x"EE", x"AA", x"EE", x"8A", x"11", x"BB", x"00", x"00", x"74", x"42", x"34", x"70", x"1A", x"3B", x"00", x"00", 
        x"77", x"55", x"56", x"75", x"15", x"D4", x"00", x"00", x"77", x"44", x"33", x"77", x"95", x"5D", x"00", x"00", 
        x"77", x"42", x"42", x"77", x"01", x"01", x"00", x"00", x"07", x"04", x"03", x"07", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"FF", x"00", x"00", x"A0", x"C0", x"A0", x"A0", x"00", x"FF", x"00", x"00", x"EE", x"A8", 
        x"A8", x"EE", x"00", x"FF", x"00", x"00", x"4E", x"2A", x"4C", x"0A", x"00", x"FF", x"00", x"00", x"77", x"45", 
        x"66", x"75", x"00", x"FF", x"00", x"00", x"77", x"55", x"77", x"54", x"00", x"FF", x"00", x"00", x"07", x"05", 
        x"07", x"04", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"4F", x"87", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FE", x"FF", x"71", x"75", x"71", 
        x"17", x"FF", x"E9", x"D0", x"FF", x"51", x"17", x"53", x"51", x"FF", x"FF", x"3F", x"FF", x"1F", x"3F", x"DF", 
        x"1F", x"FF", x"FE", x"FD", x"FF", x"11", x"55", x"31", x"57", x"FF", x"DF", x"A7", x"FF", x"FF", x"FF", x"FF", 
        x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F4", x"03", x"01", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"7D", x"3A", x"14", x"08", x"30", x"50", x"60", x"C0", x"A0", x"40", x"80", x"00", 
        x"0C", x"0A", x"06", x"03", x"1F", x"0F", x"06", x"03", x"80", x"C0", x"E0", x"20", x"FA", x"F4", x"E8", x"50", 
        x"27", x"04", x"04", x"04", x"43", x"81", x"00", x"00", x"00", x"C0", x"20", x"10", x"7F", x"3E", x"1D", x"0A", 
        x"04", x"03", x"04", x"0A", x"E8", x"D0", x"A0", x"40", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"80", x"60", x"30", x"10", x"00", x"00", x"F0", x"10", x"01", x"06", x"0C", x"08", 
        x"00", x"00", x"0F", x"08", x"20", x"20", x"20", x"E0", x"00", x"00", x"F0", x"10", x"04", x"04", x"04", x"07", 
        x"00", x"00", x"0F", x"08", x"B0", x"50", x"B0", x"60", x"C0", x"00", x"F0", x"10", x"08", x"09", x"08", x"05", 
        x"03", x"00", x"0F", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"FF", x"D0", x"10", x"10", x"D0", x"10", x"F0", x"00", x"FF", x"0B", x"0A", x"0A", x"0B", 
        x"08", x"0F", x"00", x"FF", x"50", x"90", x"90", x"50", x"10", x"F0", x"00", x"FF", x"0A", x"09", x"09", x"0A", 
        x"08", x"0F", x"00", x"FF", x"D0", x"90", x"10", x"D0", x"10", x"F0", x"00", x"FF", x"0B", x"08", x"09", x"0B", 
        x"08", x"0F", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"DE", x"5C", x"D0", 
        x"9E", x"00", x"00", x"00", x"00", x"7B", x"4A", x"4B", x"7A", x"00", x"00", x"E8", x"00", x"EF", x"08", x"E8", 
        x"EF", x"00", x"00", x"BD", x"00", x"79", x"49", x"79", x"48", x"00", x"00", x"F7", x"00", x"DE", x"48", x"48", 
        x"C8", x"00", x"00", x"BC", x"00", x"7B", x"42", x"4A", x"7B", x"00", x"00", x"97", x"00", x"D2", x"52", x"52", 
        x"DE", x"00", x"00", x"1E", x"00", x"4B", x"4A", x"7A", x"23", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"28", x"20", x"E8", x"00", x"00", x"BC", x"A4", x"BC", x"A5", x"A5", x"BD", x"00", 
        x"00", x"F7", x"84", x"E4", x"24", x"24", x"F7", x"00", x"00", x"BC", x"20", x"3C", x"24", x"3C", x"A8", x"00", 
        x"00", x"D5", x"B6", x"95", x"97", x"94", x"67", x"00", x"00", x"5E", x"52", x"DE", x"12", x"12", x"1E", x"00", 
        x"00", x"7A", x"22", x"23", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"A8", x"00", x"00", x"40", x"40", x"00", x"40", x"00", x"87", x"00", x"00", x"AF", 
        x"68", x"29", x"2F", x"00", x"9C", x"00", x"00", x"BD", x"91", x"91", x"3D", x"00", x"94", x"00", x"00", x"F4", 
        x"94", x"F7", x"92", x"00", x"52", x"00", x"00", x"D0", x"50", x"D0", x"1E", x"00", x"22", x"00", x"00", x"03", 
        x"02", x"03", x"02", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"7A", x"72", x"40", x"7A", x"00", x"00", x"00", x"00", x"EE", x"89", x"89", 
        x"EE", x"00", x"00", x"00", x"00", x"BD", x"20", x"3C", x"1D", x"00", x"00", x"00", x"00", x"97", x"92", x"92", 
        x"F2", x"00", x"00", x"00", x"00", x"9E", x"92", x"92", x"9E", x"00", x"00", x"00", x"00", x"F7", x"84", x"94", 
        x"F7", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8A", x"8A", x"AA", x"AA", 
        x"DA", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"88", x"C8", x"A8", x"98", x"88", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8E", x"8A", x"8A", x"8A", x"EE", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"88", x"EC", x"28", x"EE", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"EB", x"4A", x"4B", x"4A", x"4B", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", 
        x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", x"90", x"90", x"48", x"84", x"90", x"CD", x"FF", x"4A", 
        x"00", x"27", x"AB", x"4A", x"01", x"27", x"CD", x"4A", x"02", x"27", x"EF", x"4A", x"03", x"28", x"33", x"4A", 
        x"04", x"28", x"57", x"4A", x"05", x"28", x"11", x"17", x"8D", x"00", x"EE", x"A2", x"2C", x"28", x"3D", x"F6", 
        x"0A", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"6A", x"01", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"00", 
        x"E0", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"00", x"EE", x"17", x"AF", x"00", x"EE", x"A4", x"2C", x"28", 
        x"3D", x"F6", x"0A", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"6A", x"02", x"6E", x"00", x"8E", x"67", x"4F", 
        x"01", x"00", x"E0", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"00", x"EE", x"17", x"D1", x"00", x"EE", x"A5", 
        x"2C", x"28", x"3D", x"F6", x"0A", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"6A", x"03", x"6E", x"00", x"8E", 
        x"67", x"4F", x"01", x"00", x"E0", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"00", x"EE", x"17", x"F3", x"00", 
        x"EE", x"A6", x"2C", x"28", x"3D", x"F6", x"0A", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"6A", x"05", x"6E", 
        x"00", x"8E", x"67", x"4F", x"01", x"00", x"E0", x"6E", x"00", x"8E", x"67", x"4F", x"01", x"00", x"EE", x"18", 
        x"15", x"00", x"EE", x"A3", x"2C", x"28", x"3D", x"6A", x"04", x"29", x"A5", x"00", x"EE", x"69", x"38", x"68", 
        x"00", x"67", x"08", x"D9", x"88", x"F7", x"1E", x"79", x"F8", x"49", x"F8", x"78", x"08", x"49", x"F8", x"69", 
        x"38", x"38", x"20", x"18", x"43", x"00", x"EE", x"6E", x"00", x"8E", x"D7", x"4F", x"01", x"6C", x"01", x"6E", 
        x"56", x"8E", x"D7", x"4F", x"01", x"6C", x"02", x"6E", x"AB", x"8E", x"D7", x"4F", x"01", x"6C", x"03", x"6B", 
        x"00", x"67", x"00", x"F6", x"0A", x"46", x"0A", x"6B", x"01", x"46", x"00", x"6B", x"02", x"46", x"0B", x"6B", 
        x"03", x"4B", x"00", x"18", x"73", x"28", x"A7", x"28", x"C7", x"28", x"E7", x"29", x"67", x"35", x"01", x"18", 
        x"97", x"29", x"A5", x"70", x"01", x"29", x"A5", x"77", x"01", x"37", x"A0", x"18", x"97", x"28", x"A7", x"28", 
        x"C7", x"28", x"E7", x"29", x"67", x"00", x"EE", x"6E", x"01", x"8E", x"B7", x"4F", x"01", x"A2", x"02", x"6E", 
        x"02", x"8E", x"B7", x"4F", x"01", x"A2", x"10", x"6E", x"03", x"8E", x"B7", x"4F", x"01", x"A2", x"1E", x"69", 
        x"2C", x"68", x"0C", x"D9", x"88", x"00", x"EE", x"6E", x"01", x"8E", x"C7", x"4F", x"01", x"A2", x"02", x"6E", 
        x"02", x"8E", x"C7", x"4F", x"01", x"A2", x"10", x"6E", x"03", x"8E", x"C7", x"4F", x"01", x"A2", x"1E", x"69", 
        x"0C", x"68", x"0C", x"D9", x"88", x"00", x"EE", x"3B", x"01", x"18", x"FD", x"3C", x"01", x"18", x"F1", x"29", 
        x"53", x"3C", x"02", x"18", x"F7", x"29", x"2B", x"3C", x"03", x"18", x"FD", x"29", x"3F", x"3B", x"02", x"19", 
        x"13", x"3C", x"02", x"19", x"07", x"29", x"53", x"3C", x"03", x"19", x"0D", x"29", x"2B", x"3C", x"01", x"19", 
        x"13", x"29", x"3F", x"3B", x"03", x"19", x"29", x"3C", x"03", x"19", x"1D", x"29", x"53", x"3C", x"01", x"19", 
        x"23", x"29", x"2B", x"3C", x"02", x"19", x"29", x"29", x"3F", x"00", x"EE", x"A7", x"4A", x"69", x"01", x"68", 
        x"01", x"D9", x"85", x"A7", x"59", x"69", x"09", x"68", x"01", x"D9", x"85", x"65", x"00", x"00", x"EE", x"A7", 
        x"2C", x"69", x"01", x"68", x"01", x"D9", x"85", x"A7", x"3B", x"69", x"09", x"68", x"01", x"D9", x"85", x"65", 
        x"01", x"00", x"EE", x"A7", x"68", x"69", x"01", x"68", x"01", x"D9", x"85", x"A7", x"77", x"69", x"09", x"68", 
        x"01", x"D9", x"85", x"65", x"02", x"00", x"EE", x"35", x"00", x"19", x"7B", x"A7", x"86", x"69", x"39", x"68", 
        x"1B", x"D9", x"82", x"A7", x"88", x"69", x"03", x"68", x"1B", x"D9", x"82", x"35", x"01", x"19", x"8F", x"A7", 
        x"86", x"69", x"03", x"68", x"1B", x"D9", x"82", x"A7", x"88", x"69", x"39", x"68", x"1B", x"D9", x"82", x"35", 
        x"02", x"19", x"A3", x"A7", x"8A", x"69", x"38", x"68", x"18", x"D9", x"82", x"A7", x"88", x"69", x"03", x"68", 
        x"1C", x"D9", x"81", x"00", x"EE", x"30", x"0A", x"19", x"AD", x"71", x"01", x"60", x"00", x"31", x"0A", x"19", 
        x"B5", x"72", x"01", x"61", x"00", x"32", x"0A", x"19", x"C7", x"62", x"00", x"61", x"00", x"60", x"00", x"00", 
        x"E0", x"6A", x"05", x"27", x"8D", x"00", x"E0", x"69", x"3A", x"68", x"01", x"F0", x"29", x"D9", x"85", x"69", 
        x"35", x"68", x"01", x"F1", x"29", x"D9", x"85", x"69", x"30", x"68", x"01", x"F2", x"29", x"D9", x"85", x"00", 
        x"EE"
    );

end package;

package body rps is
end rps;